// All 12 validated RFT kernels - case statement body
// Generated from algorithms/rft/variants/operator_variants.py

            // MODE 0: RFT-GOLDEN (unitarity: 6.12e-15)
            {4'd0, 3'd0, 3'd0}: kernel_rom_out = -16'sd10528;
            {4'd0, 3'd0, 3'd1}: kernel_rom_out = 16'sd12809;
            {4'd0, 3'd0, 3'd2}: kernel_rom_out = -16'sd11788;
            {4'd0, 3'd0, 3'd3}: kernel_rom_out = -16'sd12520;
            {4'd0, 3'd0, 3'd4}: kernel_rom_out = 16'sd14036;
            {4'd0, 3'd0, 3'd5}: kernel_rom_out = -16'sd14281;
            {4'd0, 3'd0, 3'd6}: kernel_rom_out = -16'sd9488;
            {4'd0, 3'd0, 3'd7}: kernel_rom_out = -16'sd3470;
            {4'd0, 3'd1, 3'd0}: kernel_rom_out = -16'sd11613;
            {4'd0, 3'd1, 3'd1}: kernel_rom_out = 16'sd12317;
            {4'd0, 3'd1, 3'd2}: kernel_rom_out = 16'sd11248;
            {4'd0, 3'd1, 3'd3}: kernel_rom_out = -16'sd7835;
            {4'd0, 3'd1, 3'd4}: kernel_rom_out = 16'sd9793;
            {4'd0, 3'd1, 3'd5}: kernel_rom_out = 16'sd15845;
            {4'd0, 3'd1, 3'd6}: kernel_rom_out = 16'sd13399;
            {4'd0, 3'd1, 3'd7}: kernel_rom_out = 16'sd8523;
            {4'd0, 3'd2, 3'd0}: kernel_rom_out = -16'sd12087;
            {4'd0, 3'd2, 3'd1}: kernel_rom_out = -16'sd10234;
            {4'd0, 3'd2, 3'd2}: kernel_rom_out = 16'sd11353;
            {4'd0, 3'd2, 3'd3}: kernel_rom_out = -16'sd15150;
            {4'd0, 3'd2, 3'd4}: kernel_rom_out = -16'sd8738;
            {4'd0, 3'd2, 3'd5}: kernel_rom_out = 16'sd7100;
            {4'd0, 3'd2, 3'd6}: kernel_rom_out = -16'sd13620;
            {4'd0, 3'd2, 3'd7}: kernel_rom_out = -16'sd12336;
            {4'd0, 3'd3, 3'd0}: kernel_rom_out = -16'sd12043;
            {4'd0, 3'd3, 3'd1}: kernel_rom_out = -16'sd10784;
            {4'd0, 3'd3, 3'd2}: kernel_rom_out = -16'sd11936;
            {4'd0, 3'd3, 3'd3}: kernel_rom_out = -16'sd9443;
            {4'd0, 3'd3, 3'd4}: kernel_rom_out = -16'sd12944;
            {4'd0, 3'd3, 3'd5}: kernel_rom_out = -16'sd5602;
            {4'd0, 3'd3, 3'd6}: kernel_rom_out = 16'sd9043;
            {4'd0, 3'd3, 3'd7}: kernel_rom_out = 16'sd17320;
            {4'd0, 3'd4, 3'd0}: kernel_rom_out = -16'sd12043;
            {4'd0, 3'd4, 3'd1}: kernel_rom_out = 16'sd10784;
            {4'd0, 3'd4, 3'd2}: kernel_rom_out = -16'sd11936;
            {4'd0, 3'd4, 3'd3}: kernel_rom_out = 16'sd9443;
            {4'd0, 3'd4, 3'd4}: kernel_rom_out = -16'sd12944;
            {4'd0, 3'd4, 3'd5}: kernel_rom_out = 16'sd5602;
            {4'd0, 3'd4, 3'd6}: kernel_rom_out = 16'sd9043;
            {4'd0, 3'd4, 3'd7}: kernel_rom_out = -16'sd17320;
            {4'd0, 3'd5, 3'd0}: kernel_rom_out = -16'sd12087;
            {4'd0, 3'd5, 3'd1}: kernel_rom_out = 16'sd10234;
            {4'd0, 3'd5, 3'd2}: kernel_rom_out = 16'sd11353;
            {4'd0, 3'd5, 3'd3}: kernel_rom_out = 16'sd15150;
            {4'd0, 3'd5, 3'd4}: kernel_rom_out = -16'sd8738;
            {4'd0, 3'd5, 3'd5}: kernel_rom_out = -16'sd7100;
            {4'd0, 3'd5, 3'd6}: kernel_rom_out = -16'sd13620;
            {4'd0, 3'd5, 3'd7}: kernel_rom_out = 16'sd12336;
            {4'd0, 3'd6, 3'd0}: kernel_rom_out = -16'sd11613;
            {4'd0, 3'd6, 3'd1}: kernel_rom_out = -16'sd12317;
            {4'd0, 3'd6, 3'd2}: kernel_rom_out = 16'sd11248;
            {4'd0, 3'd6, 3'd3}: kernel_rom_out = 16'sd7835;
            {4'd0, 3'd6, 3'd4}: kernel_rom_out = 16'sd9793;
            {4'd0, 3'd6, 3'd5}: kernel_rom_out = -16'sd15845;
            {4'd0, 3'd6, 3'd6}: kernel_rom_out = 16'sd13399;
            {4'd0, 3'd6, 3'd7}: kernel_rom_out = -16'sd8523;
            {4'd0, 3'd7, 3'd0}: kernel_rom_out = -16'sd10528;
            {4'd0, 3'd7, 3'd1}: kernel_rom_out = -16'sd12809;
            {4'd0, 3'd7, 3'd2}: kernel_rom_out = -16'sd11788;
            {4'd0, 3'd7, 3'd3}: kernel_rom_out = 16'sd12520;
            {4'd0, 3'd7, 3'd4}: kernel_rom_out = 16'sd14036;
            {4'd0, 3'd7, 3'd5}: kernel_rom_out = 16'sd14281;
            {4'd0, 3'd7, 3'd6}: kernel_rom_out = -16'sd9488;
            {4'd0, 3'd7, 3'd7}: kernel_rom_out = 16'sd3470;

            // MODE 1: RFT-FIBONACCI (unitarity: 1.09e-13)
            {4'd1, 3'd0, 3'd0}: kernel_rom_out = 16'sd3859;
            {4'd1, 3'd0, 3'd1}: kernel_rom_out = -16'sd9620;
            {4'd1, 3'd0, 3'd2}: kernel_rom_out = 16'sd15561;
            {4'd1, 3'd0, 3'd3}: kernel_rom_out = -16'sd13362;
            {4'd1, 3'd0, 3'd4}: kernel_rom_out = 16'sd11981;
            {4'd1, 3'd0, 3'd5}: kernel_rom_out = -16'sd11555;
            {4'd1, 3'd0, 3'd6}: kernel_rom_out = 16'sd11672;
            {4'd1, 3'd0, 3'd7}: kernel_rom_out = 16'sd11499;
            {4'd1, 3'd1, 3'd0}: kernel_rom_out = 16'sd8362;
            {4'd1, 3'd1, 3'd1}: kernel_rom_out = -16'sd13352;
            {4'd1, 3'd1, 3'd2}: kernel_rom_out = 16'sd14810;
            {4'd1, 3'd1, 3'd3}: kernel_rom_out = 16'sd9564;
            {4'd1, 3'd1, 3'd4}: kernel_rom_out = -16'sd10614;
            {4'd1, 3'd1, 3'd5}: kernel_rom_out = -16'sd11499;
            {4'd1, 3'd1, 3'd6}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd1, 3'd7}: kernel_rom_out = -16'sd11613;
            {4'd1, 3'd2, 3'd0}: kernel_rom_out = 16'sd12646;
            {4'd1, 3'd2, 3'd1}: kernel_rom_out = -16'sd13286;
            {4'd1, 3'd2, 3'd2}: kernel_rom_out = -16'sd5722;
            {4'd1, 3'd2, 3'd3}: kernel_rom_out = 16'sd9516;
            {4'd1, 3'd2, 3'd4}: kernel_rom_out = 16'sd14559;
            {4'd1, 3'd2, 3'd5}: kernel_rom_out = 16'sd11614;
            {4'd1, 3'd2, 3'd6}: kernel_rom_out = -16'sd11497;
            {4'd1, 3'd2, 3'd7}: kernel_rom_out = 16'sd11613;
            {4'd1, 3'd3, 3'd0}: kernel_rom_out = 16'sd17090;
            {4'd1, 3'd3, 3'd1}: kernel_rom_out = -16'sd9460;
            {4'd1, 3'd3, 3'd2}: kernel_rom_out = -16'sd6526;
            {4'd1, 3'd3, 3'd3}: kernel_rom_out = -16'sd13276;
            {4'd1, 3'd3, 3'd4}: kernel_rom_out = -16'sd8285;
            {4'd1, 3'd3, 3'd5}: kernel_rom_out = 16'sd11671;
            {4'd1, 3'd3, 3'd6}: kernel_rom_out = 16'sd11555;
            {4'd1, 3'd3, 3'd7}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd4, 3'd0}: kernel_rom_out = 16'sd17090;
            {4'd1, 3'd4, 3'd1}: kernel_rom_out = 16'sd9460;
            {4'd1, 3'd4, 3'd2}: kernel_rom_out = -16'sd6526;
            {4'd1, 3'd4, 3'd3}: kernel_rom_out = 16'sd13276;
            {4'd1, 3'd4, 3'd4}: kernel_rom_out = -16'sd8285;
            {4'd1, 3'd4, 3'd5}: kernel_rom_out = -16'sd11671;
            {4'd1, 3'd4, 3'd6}: kernel_rom_out = 16'sd11555;
            {4'd1, 3'd4, 3'd7}: kernel_rom_out = 16'sd11614;
            {4'd1, 3'd5, 3'd0}: kernel_rom_out = 16'sd12646;
            {4'd1, 3'd5, 3'd1}: kernel_rom_out = 16'sd13286;
            {4'd1, 3'd5, 3'd2}: kernel_rom_out = -16'sd5722;
            {4'd1, 3'd5, 3'd3}: kernel_rom_out = -16'sd9516;
            {4'd1, 3'd5, 3'd4}: kernel_rom_out = 16'sd14559;
            {4'd1, 3'd5, 3'd5}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd5, 3'd6}: kernel_rom_out = -16'sd11497;
            {4'd1, 3'd5, 3'd7}: kernel_rom_out = -16'sd11613;
            {4'd1, 3'd6, 3'd0}: kernel_rom_out = 16'sd8362;
            {4'd1, 3'd6, 3'd1}: kernel_rom_out = 16'sd13352;
            {4'd1, 3'd6, 3'd2}: kernel_rom_out = 16'sd14810;
            {4'd1, 3'd6, 3'd3}: kernel_rom_out = -16'sd9564;
            {4'd1, 3'd6, 3'd4}: kernel_rom_out = -16'sd10614;
            {4'd1, 3'd6, 3'd5}: kernel_rom_out = 16'sd11499;
            {4'd1, 3'd6, 3'd6}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd6, 3'd7}: kernel_rom_out = 16'sd11613;
            {4'd1, 3'd7, 3'd0}: kernel_rom_out = 16'sd3859;
            {4'd1, 3'd7, 3'd1}: kernel_rom_out = 16'sd9620;
            {4'd1, 3'd7, 3'd2}: kernel_rom_out = 16'sd15561;
            {4'd1, 3'd7, 3'd3}: kernel_rom_out = 16'sd13362;
            {4'd1, 3'd7, 3'd4}: kernel_rom_out = 16'sd11981;
            {4'd1, 3'd7, 3'd5}: kernel_rom_out = 16'sd11555;
            {4'd1, 3'd7, 3'd6}: kernel_rom_out = 16'sd11672;
            {4'd1, 3'd7, 3'd7}: kernel_rom_out = -16'sd11499;

            // MODE 2: RFT-HARMONIC (unitarity: 1.96e-15)
            {4'd2, 3'd0, 3'd0}: kernel_rom_out = 16'sd11505;
            {4'd2, 3'd0, 3'd1}: kernel_rom_out = -16'sd11573;
            {4'd2, 3'd0, 3'd2}: kernel_rom_out = 16'sd14539;
            {4'd2, 3'd0, 3'd3}: kernel_rom_out = 16'sd16484;
            {4'd2, 3'd0, 3'd4}: kernel_rom_out = 16'sd8842;
            {4'd2, 3'd0, 3'd5}: kernel_rom_out = -16'sd13592;
            {4'd2, 3'd0, 3'd6}: kernel_rom_out = 16'sd2596;
            {4'd2, 3'd0, 3'd7}: kernel_rom_out = 16'sd7386;
            {4'd2, 3'd1, 3'd0}: kernel_rom_out = -16'sd11549;
            {4'd2, 3'd1, 3'd1}: kernel_rom_out = -16'sd11481;
            {4'd2, 3'd1, 3'd2}: kernel_rom_out = -16'sd15661;
            {4'd2, 3'd1, 3'd3}: kernel_rom_out = 16'sd13444;
            {4'd2, 3'd1, 3'd4}: kernel_rom_out = -16'sd14106;
            {4'd2, 3'd1, 3'd5}: kernel_rom_out = -16'sd8723;
            {4'd2, 3'd1, 3'd6}: kernel_rom_out = -16'sd9147;
            {4'd2, 3'd1, 3'd7}: kernel_rom_out = 16'sd4871;
            {4'd2, 3'd2, 3'd0}: kernel_rom_out = 16'sd11635;
            {4'd2, 3'd2, 3'd1}: kernel_rom_out = -16'sd11657;
            {4'd2, 3'd2, 3'd2}: kernel_rom_out = 16'sd6800;
            {4'd2, 3'd2, 3'd3}: kernel_rom_out = 16'sd4852;
            {4'd2, 3'd2, 3'd4}: kernel_rom_out = -16'sd10542;
            {4'd2, 3'd2, 3'd5}: kernel_rom_out = 16'sd15032;
            {4'd2, 3'd2, 3'd6}: kernel_rom_out = -16'sd11345;
            {4'd2, 3'd2, 3'd7}: kernel_rom_out = -16'sd16334;
            {4'd2, 3'd3, 3'd0}: kernel_rom_out = -16'sd11649;
            {4'd2, 3'd3, 3'd1}: kernel_rom_out = -16'sd11626;
            {4'd2, 3'd3, 3'd2}: kernel_rom_out = -16'sd5826;
            {4'd2, 3'd3, 3'd3}: kernel_rom_out = 16'sd7797;
            {4'd2, 3'd3, 3'd4}: kernel_rom_out = 16'sd12188;
            {4'd2, 3'd3, 3'd5}: kernel_rom_out = 16'sd7072;
            {4'd2, 3'd3, 3'd6}: kernel_rom_out = 16'sd17824;
            {4'd2, 3'd3, 3'd7}: kernel_rom_out = -16'sd13848;
            {4'd2, 3'd4, 3'd0}: kernel_rom_out = 16'sd11649;
            {4'd2, 3'd4, 3'd1}: kernel_rom_out = -16'sd11626;
            {4'd2, 3'd4, 3'd2}: kernel_rom_out = -16'sd5826;
            {4'd2, 3'd4, 3'd3}: kernel_rom_out = -16'sd7797;
            {4'd2, 3'd4, 3'd4}: kernel_rom_out = -16'sd12188;
            {4'd2, 3'd4, 3'd5}: kernel_rom_out = 16'sd7072;
            {4'd2, 3'd4, 3'd6}: kernel_rom_out = 16'sd17824;
            {4'd2, 3'd4, 3'd7}: kernel_rom_out = 16'sd13848;
            {4'd2, 3'd5, 3'd0}: kernel_rom_out = -16'sd11635;
            {4'd2, 3'd5, 3'd1}: kernel_rom_out = -16'sd11657;
            {4'd2, 3'd5, 3'd2}: kernel_rom_out = 16'sd6800;
            {4'd2, 3'd5, 3'd3}: kernel_rom_out = -16'sd4852;
            {4'd2, 3'd5, 3'd4}: kernel_rom_out = 16'sd10542;
            {4'd2, 3'd5, 3'd5}: kernel_rom_out = 16'sd15032;
            {4'd2, 3'd5, 3'd6}: kernel_rom_out = -16'sd11345;
            {4'd2, 3'd5, 3'd7}: kernel_rom_out = 16'sd16334;
            {4'd2, 3'd6, 3'd0}: kernel_rom_out = 16'sd11549;
            {4'd2, 3'd6, 3'd1}: kernel_rom_out = -16'sd11481;
            {4'd2, 3'd6, 3'd2}: kernel_rom_out = -16'sd15661;
            {4'd2, 3'd6, 3'd3}: kernel_rom_out = -16'sd13444;
            {4'd2, 3'd6, 3'd4}: kernel_rom_out = 16'sd14106;
            {4'd2, 3'd6, 3'd5}: kernel_rom_out = -16'sd8723;
            {4'd2, 3'd6, 3'd6}: kernel_rom_out = -16'sd9147;
            {4'd2, 3'd6, 3'd7}: kernel_rom_out = -16'sd4871;
            {4'd2, 3'd7, 3'd0}: kernel_rom_out = -16'sd11505;
            {4'd2, 3'd7, 3'd1}: kernel_rom_out = -16'sd11573;
            {4'd2, 3'd7, 3'd2}: kernel_rom_out = 16'sd14539;
            {4'd2, 3'd7, 3'd3}: kernel_rom_out = -16'sd16484;
            {4'd2, 3'd7, 3'd4}: kernel_rom_out = -16'sd8842;
            {4'd2, 3'd7, 3'd5}: kernel_rom_out = -16'sd13592;
            {4'd2, 3'd7, 3'd6}: kernel_rom_out = 16'sd2596;
            {4'd2, 3'd7, 3'd7}: kernel_rom_out = -16'sd7386;

            // MODE 3: RFT-GEOMETRIC (unitarity: 3.58e-15)
            {4'd3, 3'd0, 3'd0}: kernel_rom_out = -16'sd13692;
            {4'd3, 3'd0, 3'd1}: kernel_rom_out = 16'sd663;
            {4'd3, 3'd0, 3'd2}: kernel_rom_out = 16'sd20505;
            {4'd3, 3'd0, 3'd3}: kernel_rom_out = -16'sd9236;
            {4'd3, 3'd0, 3'd4}: kernel_rom_out = -16'sd9709;
            {4'd3, 3'd0, 3'd5}: kernel_rom_out = -16'sd3379;
            {4'd3, 3'd0, 3'd6}: kernel_rom_out = 16'sd15895;
            {4'd3, 3'd0, 3'd7}: kernel_rom_out = -16'sd4653;
            {4'd3, 3'd1, 3'd0}: kernel_rom_out = -16'sd10201;
            {4'd3, 3'd1, 3'd1}: kernel_rom_out = 16'sd13503;
            {4'd3, 3'd1, 3'd2}: kernel_rom_out = 16'sd8329;
            {4'd3, 3'd1, 3'd3}: kernel_rom_out = 16'sd4498;
            {4'd3, 3'd1, 3'd4}: kernel_rom_out = 16'sd13956;
            {4'd3, 3'd1, 3'd5}: kernel_rom_out = 16'sd20225;
            {4'd3, 3'd1, 3'd6}: kernel_rom_out = -16'sd1874;
            {4'd3, 3'd1, 3'd7}: kernel_rom_out = 16'sd9506;
            {4'd3, 3'd2, 3'd0}: kernel_rom_out = 16'sd4467;
            {4'd3, 3'd2, 3'd1}: kernel_rom_out = 16'sd17252;
            {4'd3, 3'd2, 3'd2}: kernel_rom_out = -16'sd5562;
            {4'd3, 3'd2, 3'd3}: kernel_rom_out = 16'sd17817;
            {4'd3, 3'd2, 3'd4}: kernel_rom_out = -16'sd3910;
            {4'd3, 3'd2, 3'd5}: kernel_rom_out = -16'sd401;
            {4'd3, 3'd2, 3'd6}: kernel_rom_out = 16'sd14116;
            {4'd3, 3'd2, 3'd7}: kernel_rom_out = -16'sd13892;
            {4'd3, 3'd3, 3'd0}: kernel_rom_out = 16'sd15012;
            {4'd3, 3'd3, 3'd1}: kernel_rom_out = 16'sd7512;
            {4'd3, 3'd3, 3'd2}: kernel_rom_out = -16'sd4007;
            {4'd3, 3'd3, 3'd3}: kernel_rom_out = -16'sd10670;
            {4'd3, 3'd3, 3'd4}: kernel_rom_out = -16'sd15248;
            {4'd3, 3'd3, 3'd5}: kernel_rom_out = 16'sd10781;
            {4'd3, 3'd3, 3'd6}: kernel_rom_out = 16'sd9023;
            {4'd3, 3'd3, 3'd7}: kernel_rom_out = 16'sd15226;
            {4'd3, 3'd4, 3'd0}: kernel_rom_out = 16'sd15012;
            {4'd3, 3'd4, 3'd1}: kernel_rom_out = -16'sd7512;
            {4'd3, 3'd4, 3'd2}: kernel_rom_out = 16'sd4007;
            {4'd3, 3'd4, 3'd3}: kernel_rom_out = -16'sd10670;
            {4'd3, 3'd4, 3'd4}: kernel_rom_out = 16'sd15248;
            {4'd3, 3'd4, 3'd5}: kernel_rom_out = 16'sd10781;
            {4'd3, 3'd4, 3'd6}: kernel_rom_out = 16'sd9023;
            {4'd3, 3'd4, 3'd7}: kernel_rom_out = -16'sd15226;
            {4'd3, 3'd5, 3'd0}: kernel_rom_out = 16'sd4467;
            {4'd3, 3'd5, 3'd1}: kernel_rom_out = -16'sd17252;
            {4'd3, 3'd5, 3'd2}: kernel_rom_out = 16'sd5562;
            {4'd3, 3'd5, 3'd3}: kernel_rom_out = 16'sd17817;
            {4'd3, 3'd5, 3'd4}: kernel_rom_out = 16'sd3910;
            {4'd3, 3'd5, 3'd5}: kernel_rom_out = -16'sd401;
            {4'd3, 3'd5, 3'd6}: kernel_rom_out = 16'sd14116;
            {4'd3, 3'd5, 3'd7}: kernel_rom_out = 16'sd13892;
            {4'd3, 3'd6, 3'd0}: kernel_rom_out = -16'sd10201;
            {4'd3, 3'd6, 3'd1}: kernel_rom_out = -16'sd13503;
            {4'd3, 3'd6, 3'd2}: kernel_rom_out = -16'sd8329;
            {4'd3, 3'd6, 3'd3}: kernel_rom_out = 16'sd4498;
            {4'd3, 3'd6, 3'd4}: kernel_rom_out = -16'sd13956;
            {4'd3, 3'd6, 3'd5}: kernel_rom_out = 16'sd20225;
            {4'd3, 3'd6, 3'd6}: kernel_rom_out = -16'sd1874;
            {4'd3, 3'd6, 3'd7}: kernel_rom_out = -16'sd9506;
            {4'd3, 3'd7, 3'd0}: kernel_rom_out = -16'sd13692;
            {4'd3, 3'd7, 3'd1}: kernel_rom_out = -16'sd663;
            {4'd3, 3'd7, 3'd2}: kernel_rom_out = -16'sd20505;
            {4'd3, 3'd7, 3'd3}: kernel_rom_out = -16'sd9236;
            {4'd3, 3'd7, 3'd4}: kernel_rom_out = 16'sd9709;
            {4'd3, 3'd7, 3'd5}: kernel_rom_out = -16'sd3379;
            {4'd3, 3'd7, 3'd6}: kernel_rom_out = 16'sd15895;
            {4'd3, 3'd7, 3'd7}: kernel_rom_out = 16'sd4653;

            // MODE 4: RFT-BEATING (unitarity: 3.09e-15)
            {4'd4, 3'd0, 3'd0}: kernel_rom_out = -16'sd11094;
            {4'd4, 3'd0, 3'd1}: kernel_rom_out = 16'sd15417;
            {4'd4, 3'd0, 3'd2}: kernel_rom_out = 16'sd5892;
            {4'd4, 3'd0, 3'd3}: kernel_rom_out = -16'sd12981;
            {4'd4, 3'd0, 3'd4}: kernel_rom_out = 16'sd18457;
            {4'd4, 3'd0, 3'd5}: kernel_rom_out = -16'sd6279;
            {4'd4, 3'd0, 3'd6}: kernel_rom_out = 16'sd6194;
            {4'd4, 3'd0, 3'd7}: kernel_rom_out = -16'sd9551;
            {4'd4, 3'd1, 3'd0}: kernel_rom_out = -16'sd12220;
            {4'd4, 3'd1, 3'd1}: kernel_rom_out = -16'sd6858;
            {4'd4, 3'd1, 3'd2}: kernel_rom_out = -16'sd14172;
            {4'd4, 3'd1, 3'd3}: kernel_rom_out = -16'sd16386;
            {4'd4, 3'd1, 3'd4}: kernel_rom_out = -16'sd6798;
            {4'd4, 3'd1, 3'd5}: kernel_rom_out = 16'sd14804;
            {4'd4, 3'd1, 3'd6}: kernel_rom_out = 16'sd11852;
            {4'd4, 3'd1, 3'd7}: kernel_rom_out = 16'sd1466;
            {4'd4, 3'd2, 3'd0}: kernel_rom_out = -16'sd10860;
            {4'd4, 3'd2, 3'd1}: kernel_rom_out = -16'sd5461;
            {4'd4, 3'd2, 3'd2}: kernel_rom_out = 16'sd16367;
            {4'd4, 3'd2, 3'd3}: kernel_rom_out = -16'sd9717;
            {4'd4, 3'd2, 3'd4}: kernel_rom_out = -16'sd12212;
            {4'd4, 3'd2, 3'd5}: kernel_rom_out = -16'sd14677;
            {4'd4, 3'd2, 3'd6}: kernel_rom_out = 16'sd1369;
            {4'd4, 3'd2, 3'd7}: kernel_rom_out = 16'sd14042;
            {4'd4, 3'd3, 3'd0}: kernel_rom_out = -16'sd12104;
            {4'd4, 3'd3, 3'd1}: kernel_rom_out = 16'sd14909;
            {4'd4, 3'd3, 3'd2}: kernel_rom_out = -16'sd5778;
            {4'd4, 3'd3, 3'd3}: kernel_rom_out = 16'sd2326;
            {4'd4, 3'd3, 3'd4}: kernel_rom_out = 16'sd903;
            {4'd4, 3'd3, 3'd5}: kernel_rom_out = 16'sd7927;
            {4'd4, 3'd3, 3'd6}: kernel_rom_out = -16'sd18871;
            {4'd4, 3'd3, 3'd7}: kernel_rom_out = 16'sd15694;
            {4'd4, 3'd4, 3'd0}: kernel_rom_out = -16'sd12104;
            {4'd4, 3'd4, 3'd1}: kernel_rom_out = -16'sd14909;
            {4'd4, 3'd4, 3'd2}: kernel_rom_out = -16'sd5778;
            {4'd4, 3'd4, 3'd3}: kernel_rom_out = -16'sd2326;
            {4'd4, 3'd4, 3'd4}: kernel_rom_out = 16'sd903;
            {4'd4, 3'd4, 3'd5}: kernel_rom_out = -16'sd7927;
            {4'd4, 3'd4, 3'd6}: kernel_rom_out = -16'sd18871;
            {4'd4, 3'd4, 3'd7}: kernel_rom_out = -16'sd15694;
            {4'd4, 3'd5, 3'd0}: kernel_rom_out = -16'sd10860;
            {4'd4, 3'd5, 3'd1}: kernel_rom_out = 16'sd5461;
            {4'd4, 3'd5, 3'd2}: kernel_rom_out = 16'sd16367;
            {4'd4, 3'd5, 3'd3}: kernel_rom_out = 16'sd9717;
            {4'd4, 3'd5, 3'd4}: kernel_rom_out = -16'sd12212;
            {4'd4, 3'd5, 3'd5}: kernel_rom_out = 16'sd14677;
            {4'd4, 3'd5, 3'd6}: kernel_rom_out = 16'sd1369;
            {4'd4, 3'd5, 3'd7}: kernel_rom_out = -16'sd14042;
            {4'd4, 3'd6, 3'd0}: kernel_rom_out = -16'sd12220;
            {4'd4, 3'd6, 3'd1}: kernel_rom_out = 16'sd6858;
            {4'd4, 3'd6, 3'd2}: kernel_rom_out = -16'sd14172;
            {4'd4, 3'd6, 3'd3}: kernel_rom_out = 16'sd16386;
            {4'd4, 3'd6, 3'd4}: kernel_rom_out = -16'sd6798;
            {4'd4, 3'd6, 3'd5}: kernel_rom_out = -16'sd14804;
            {4'd4, 3'd6, 3'd6}: kernel_rom_out = 16'sd11852;
            {4'd4, 3'd6, 3'd7}: kernel_rom_out = -16'sd1466;
            {4'd4, 3'd7, 3'd0}: kernel_rom_out = -16'sd11094;
            {4'd4, 3'd7, 3'd1}: kernel_rom_out = -16'sd15417;
            {4'd4, 3'd7, 3'd2}: kernel_rom_out = 16'sd5892;
            {4'd4, 3'd7, 3'd3}: kernel_rom_out = 16'sd12981;
            {4'd4, 3'd7, 3'd4}: kernel_rom_out = 16'sd18457;
            {4'd4, 3'd7, 3'd5}: kernel_rom_out = 16'sd6279;
            {4'd4, 3'd7, 3'd6}: kernel_rom_out = 16'sd6194;
            {4'd4, 3'd7, 3'd7}: kernel_rom_out = 16'sd9551;

            // MODE 5: RFT-PHYLLOTAXIS (unitarity: 4.38e-15)
            {4'd5, 3'd0, 3'd0}: kernel_rom_out = 16'sd9597;
            {4'd5, 3'd0, 3'd1}: kernel_rom_out = 16'sd15505;
            {4'd5, 3'd0, 3'd2}: kernel_rom_out = -16'sd9608;
            {4'd5, 3'd0, 3'd3}: kernel_rom_out = 16'sd5574;
            {4'd5, 3'd0, 3'd4}: kernel_rom_out = 16'sd13824;
            {4'd5, 3'd0, 3'd5}: kernel_rom_out = -16'sd3604;
            {4'd5, 3'd0, 3'd6}: kernel_rom_out = 16'sd16222;
            {4'd5, 3'd0, 3'd7}: kernel_rom_out = -16'sd12268;
            {4'd5, 3'd1, 3'd0}: kernel_rom_out = -16'sd16171;
            {4'd5, 3'd1, 3'd1}: kernel_rom_out = -16'sd1835;
            {4'd5, 3'd1, 3'd2}: kernel_rom_out = 16'sd248;
            {4'd5, 3'd1, 3'd3}: kernel_rom_out = 16'sd12282;
            {4'd5, 3'd1, 3'd4}: kernel_rom_out = 16'sd7890;
            {4'd5, 3'd1, 3'd5}: kernel_rom_out = 16'sd21706;
            {4'd5, 3'd1, 3'd6}: kernel_rom_out = -16'sd2818;
            {4'd5, 3'd1, 3'd7}: kernel_rom_out = -16'sd10796;
            {4'd5, 3'd2, 3'd0}: kernel_rom_out = 16'sd12685;
            {4'd5, 3'd2, 3'd1}: kernel_rom_out = -16'sd11019;
            {4'd5, 3'd2, 3'd2}: kernel_rom_out = 16'sd9066;
            {4'd5, 3'd2, 3'd3}: kernel_rom_out = 16'sd4638;
            {4'd5, 3'd2, 3'd4}: kernel_rom_out = 16'sd16799;
            {4'd5, 3'd2, 3'd5}: kernel_rom_out = -16'sd7142;
            {4'd5, 3'd2, 3'd6}: kernel_rom_out = -16'sd16266;
            {4'd5, 3'd2, 3'd7}: kernel_rom_out = -16'sd9477;
            {4'd5, 3'd3, 3'd0}: kernel_rom_out = -16'sd4725;
            {4'd5, 3'd3, 3'd1}: kernel_rom_out = 16'sd13100;
            {4'd5, 3'd3, 3'd2}: kernel_rom_out = 16'sd19033;
            {4'd5, 3'd3, 3'd3}: kernel_rom_out = -16'sd18259;
            {4'd5, 3'd3, 3'd4}: kernel_rom_out = -16'sd1126;
            {4'd5, 3'd3, 3'd5}: kernel_rom_out = 16'sd1299;
            {4'd5, 3'd3, 3'd6}: kernel_rom_out = -16'sd1075;
            {4'd5, 3'd3, 3'd7}: kernel_rom_out = -16'sd13415;
            {4'd5, 3'd4, 3'd0}: kernel_rom_out = -16'sd4725;
            {4'd5, 3'd4, 3'd1}: kernel_rom_out = -16'sd13100;
            {4'd5, 3'd4, 3'd2}: kernel_rom_out = -16'sd19033;
            {4'd5, 3'd4, 3'd3}: kernel_rom_out = -16'sd18259;
            {4'd5, 3'd4, 3'd4}: kernel_rom_out = 16'sd1126;
            {4'd5, 3'd4, 3'd5}: kernel_rom_out = -16'sd1299;
            {4'd5, 3'd4, 3'd6}: kernel_rom_out = -16'sd1075;
            {4'd5, 3'd4, 3'd7}: kernel_rom_out = -16'sd13415;
            {4'd5, 3'd5, 3'd0}: kernel_rom_out = 16'sd12685;
            {4'd5, 3'd5, 3'd1}: kernel_rom_out = 16'sd11019;
            {4'd5, 3'd5, 3'd2}: kernel_rom_out = -16'sd9066;
            {4'd5, 3'd5, 3'd3}: kernel_rom_out = 16'sd4638;
            {4'd5, 3'd5, 3'd4}: kernel_rom_out = -16'sd16799;
            {4'd5, 3'd5, 3'd5}: kernel_rom_out = 16'sd7142;
            {4'd5, 3'd5, 3'd6}: kernel_rom_out = -16'sd16266;
            {4'd5, 3'd5, 3'd7}: kernel_rom_out = -16'sd9477;
            {4'd5, 3'd6, 3'd0}: kernel_rom_out = -16'sd16171;
            {4'd5, 3'd6, 3'd1}: kernel_rom_out = 16'sd1835;
            {4'd5, 3'd6, 3'd2}: kernel_rom_out = -16'sd248;
            {4'd5, 3'd6, 3'd3}: kernel_rom_out = 16'sd12282;
            {4'd5, 3'd6, 3'd4}: kernel_rom_out = -16'sd7890;
            {4'd5, 3'd6, 3'd5}: kernel_rom_out = -16'sd21706;
            {4'd5, 3'd6, 3'd6}: kernel_rom_out = -16'sd2818;
            {4'd5, 3'd6, 3'd7}: kernel_rom_out = -16'sd10796;
            {4'd5, 3'd7, 3'd0}: kernel_rom_out = 16'sd9597;
            {4'd5, 3'd7, 3'd1}: kernel_rom_out = -16'sd15505;
            {4'd5, 3'd7, 3'd2}: kernel_rom_out = 16'sd9608;
            {4'd5, 3'd7, 3'd3}: kernel_rom_out = 16'sd5574;
            {4'd5, 3'd7, 3'd4}: kernel_rom_out = -16'sd13824;
            {4'd5, 3'd7, 3'd5}: kernel_rom_out = 16'sd3604;
            {4'd5, 3'd7, 3'd6}: kernel_rom_out = 16'sd16222;
            {4'd5, 3'd7, 3'd7}: kernel_rom_out = -16'sd12268;

            // MODE 6: RFT-CASCADE (unitarity: 1.51e-15)
            {4'd6, 3'd0, 3'd0}: kernel_rom_out = -16'sd9727;
            {4'd6, 3'd0, 3'd1}: kernel_rom_out = 16'sd15910;
            {4'd6, 3'd0, 3'd2}: kernel_rom_out = 16'sd14164;
            {4'd6, 3'd0, 3'd3}: kernel_rom_out = -16'sd2527;
            {4'd6, 3'd0, 3'd4}: kernel_rom_out = 16'sd15410;
            {4'd6, 3'd0, 3'd5}: kernel_rom_out = -16'sd4311;
            {4'd6, 3'd0, 3'd6}: kernel_rom_out = 16'sd2029;
            {4'd6, 3'd0, 3'd7}: kernel_rom_out = 16'sd16085;
            {4'd6, 3'd1, 3'd0}: kernel_rom_out = -16'sd10888;
            {4'd6, 3'd1, 3'd1}: kernel_rom_out = 16'sd16012;
            {4'd6, 3'd1, 3'd2}: kernel_rom_out = -16'sd12647;
            {4'd6, 3'd1, 3'd3}: kernel_rom_out = -16'sd3171;
            {4'd6, 3'd1, 3'd4}: kernel_rom_out = 16'sd2664;
            {4'd6, 3'd1, 3'd5}: kernel_rom_out = 16'sd8553;
            {4'd6, 3'd1, 3'd6}: kernel_rom_out = 16'sd15851;
            {4'd6, 3'd1, 3'd7}: kernel_rom_out = -16'sd14044;
            {4'd6, 3'd2, 3'd0}: kernel_rom_out = -16'sd12549;
            {4'd6, 3'd2, 3'd1}: kernel_rom_out = -16'sd1629;
            {4'd6, 3'd2, 3'd2}: kernel_rom_out = -16'sd9517;
            {4'd6, 3'd2, 3'd3}: kernel_rom_out = -16'sd19434;
            {4'd6, 3'd2, 3'd4}: kernel_rom_out = 16'sd3029;
            {4'd6, 3'd2, 3'd5}: kernel_rom_out = -16'sd11648;
            {4'd6, 3'd2, 3'd6}: kernel_rom_out = -16'sd16722;
            {4'd6, 3'd2, 3'd7}: kernel_rom_out = -16'sd4564;
            {4'd6, 3'd3, 3'd0}: kernel_rom_out = -16'sd12892;
            {4'd6, 3'd3, 3'd1}: kernel_rom_out = -16'sd4965;
            {4'd6, 3'd3, 3'd2}: kernel_rom_out = 16'sd9257;
            {4'd6, 3'd3, 3'd3}: kernel_rom_out = -16'sd11946;
            {4'd6, 3'd3, 3'd4}: kernel_rom_out = -16'sd16825;
            {4'd6, 3'd3, 3'd5}: kernel_rom_out = 16'sd17590;
            {4'd6, 3'd3, 3'd6}: kernel_rom_out = 16'sd1358;
            {4'd6, 3'd3, 3'd7}: kernel_rom_out = 16'sd7749;
            {4'd6, 3'd4, 3'd0}: kernel_rom_out = -16'sd12892;
            {4'd6, 3'd4, 3'd1}: kernel_rom_out = 16'sd4965;
            {4'd6, 3'd4, 3'd2}: kernel_rom_out = 16'sd9257;
            {4'd6, 3'd4, 3'd3}: kernel_rom_out = 16'sd11946;
            {4'd6, 3'd4, 3'd4}: kernel_rom_out = -16'sd16825;
            {4'd6, 3'd4, 3'd5}: kernel_rom_out = -16'sd17590;
            {4'd6, 3'd4, 3'd6}: kernel_rom_out = 16'sd1358;
            {4'd6, 3'd4, 3'd7}: kernel_rom_out = -16'sd7749;
            {4'd6, 3'd5, 3'd0}: kernel_rom_out = -16'sd12549;
            {4'd6, 3'd5, 3'd1}: kernel_rom_out = 16'sd1629;
            {4'd6, 3'd5, 3'd2}: kernel_rom_out = -16'sd9517;
            {4'd6, 3'd5, 3'd3}: kernel_rom_out = 16'sd19434;
            {4'd6, 3'd5, 3'd4}: kernel_rom_out = 16'sd3029;
            {4'd6, 3'd5, 3'd5}: kernel_rom_out = 16'sd11648;
            {4'd6, 3'd5, 3'd6}: kernel_rom_out = -16'sd16722;
            {4'd6, 3'd5, 3'd7}: kernel_rom_out = 16'sd4564;
            {4'd6, 3'd6, 3'd0}: kernel_rom_out = -16'sd10888;
            {4'd6, 3'd6, 3'd1}: kernel_rom_out = -16'sd16012;
            {4'd6, 3'd6, 3'd2}: kernel_rom_out = -16'sd12647;
            {4'd6, 3'd6, 3'd3}: kernel_rom_out = 16'sd3171;
            {4'd6, 3'd6, 3'd4}: kernel_rom_out = 16'sd2664;
            {4'd6, 3'd6, 3'd5}: kernel_rom_out = -16'sd8553;
            {4'd6, 3'd6, 3'd6}: kernel_rom_out = 16'sd15851;
            {4'd6, 3'd6, 3'd7}: kernel_rom_out = 16'sd14044;
            {4'd6, 3'd7, 3'd0}: kernel_rom_out = -16'sd9727;
            {4'd6, 3'd7, 3'd1}: kernel_rom_out = -16'sd15910;
            {4'd6, 3'd7, 3'd2}: kernel_rom_out = 16'sd14164;
            {4'd6, 3'd7, 3'd3}: kernel_rom_out = 16'sd2527;
            {4'd6, 3'd7, 3'd4}: kernel_rom_out = 16'sd15410;
            {4'd6, 3'd7, 3'd5}: kernel_rom_out = 16'sd4311;
            {4'd6, 3'd7, 3'd6}: kernel_rom_out = 16'sd2029;
            {4'd6, 3'd7, 3'd7}: kernel_rom_out = -16'sd16085;

            // MODE 7: RFT-HYBRID_DCT (unitarity: 1.12e-15)
            {4'd7, 3'd0, 3'd0}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd1}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd2}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd3}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd4}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd5}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd6}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd7}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd1, 3'd0}: kernel_rom_out = -16'sd16069;
            {4'd7, 3'd1, 3'd1}: kernel_rom_out = -16'sd13622;
            {4'd7, 3'd1, 3'd2}: kernel_rom_out = -16'sd9102;
            {4'd7, 3'd1, 3'd3}: kernel_rom_out = -16'sd3196;
            {4'd7, 3'd1, 3'd4}: kernel_rom_out = 16'sd3196;
            {4'd7, 3'd1, 3'd5}: kernel_rom_out = 16'sd9102;
            {4'd7, 3'd1, 3'd6}: kernel_rom_out = 16'sd13622;
            {4'd7, 3'd1, 3'd7}: kernel_rom_out = 16'sd16069;
            {4'd7, 3'd2, 3'd0}: kernel_rom_out = 16'sd15136;
            {4'd7, 3'd2, 3'd1}: kernel_rom_out = 16'sd6269;
            {4'd7, 3'd2, 3'd2}: kernel_rom_out = -16'sd6269;
            {4'd7, 3'd2, 3'd3}: kernel_rom_out = -16'sd15136;
            {4'd7, 3'd2, 3'd4}: kernel_rom_out = -16'sd15136;
            {4'd7, 3'd2, 3'd5}: kernel_rom_out = -16'sd6269;
            {4'd7, 3'd2, 3'd6}: kernel_rom_out = 16'sd6269;
            {4'd7, 3'd2, 3'd7}: kernel_rom_out = 16'sd15136;
            {4'd7, 3'd3, 3'd0}: kernel_rom_out = 16'sd13622;
            {4'd7, 3'd3, 3'd1}: kernel_rom_out = -16'sd3196;
            {4'd7, 3'd3, 3'd2}: kernel_rom_out = -16'sd16069;
            {4'd7, 3'd3, 3'd3}: kernel_rom_out = -16'sd9102;
            {4'd7, 3'd3, 3'd4}: kernel_rom_out = 16'sd9102;
            {4'd7, 3'd3, 3'd5}: kernel_rom_out = 16'sd16069;
            {4'd7, 3'd3, 3'd6}: kernel_rom_out = 16'sd3196;
            {4'd7, 3'd3, 3'd7}: kernel_rom_out = -16'sd13622;
            {4'd7, 3'd4, 3'd0}: kernel_rom_out = -16'sd9051;
            {4'd7, 3'd4, 3'd1}: kernel_rom_out = 16'sd15560;
            {4'd7, 3'd4, 3'd2}: kernel_rom_out = -16'sd9371;
            {4'd7, 3'd4, 3'd3}: kernel_rom_out = 16'sd10393;
            {4'd7, 3'd4, 3'd4}: kernel_rom_out = -16'sd15759;
            {4'd7, 3'd4, 3'd5}: kernel_rom_out = 16'sd4982;
            {4'd7, 3'd4, 3'd6}: kernel_rom_out = 16'sd13356;
            {4'd7, 3'd4, 3'd7}: kernel_rom_out = -16'sd10111;
            {4'd7, 3'd5, 3'd0}: kernel_rom_out = 16'sd2248;
            {4'd7, 3'd5, 3'd1}: kernel_rom_out = -16'sd7751;
            {4'd7, 3'd5, 3'd2}: kernel_rom_out = 16'sd10583;
            {4'd7, 3'd5, 3'd3}: kernel_rom_out = -16'sd6173;
            {4'd7, 3'd5, 3'd4}: kernel_rom_out = 16'sd3647;
            {4'd7, 3'd5, 3'd5}: kernel_rom_out = -16'sd13262;
            {4'd7, 3'd5, 3'd6}: kernel_rom_out = 16'sd22846;
            {4'd7, 3'd5, 3'd7}: kernel_rom_out = -16'sd12137;
            {4'd7, 3'd6, 3'd0}: kernel_rom_out = -16'sd7156;
            {4'd7, 3'd6, 3'd1}: kernel_rom_out = 16'sd3009;
            {4'd7, 3'd6, 3'd2}: kernel_rom_out = 16'sd18306;
            {4'd7, 3'd6, 3'd3}: kernel_rom_out = -16'sd16873;
            {4'd7, 3'd6, 3'd4}: kernel_rom_out = -16'sd8604;
            {4'd7, 3'd6, 3'd5}: kernel_rom_out = 16'sd17310;
            {4'd7, 3'd6, 3'd6}: kernel_rom_out = -16'sd2008;
            {4'd7, 3'd6, 3'd7}: kernel_rom_out = -16'sd3983;
            {4'd7, 3'd7, 3'd0}: kernel_rom_out = -16'sd11331;
            {4'd7, 3'd7, 3'd1}: kernel_rom_out = 16'sd19827;
            {4'd7, 3'd7, 3'd2}: kernel_rom_out = -16'sd4917;
            {4'd7, 3'd7, 3'd3}: kernel_rom_out = -16'sd13655;
            {4'd7, 3'd7, 3'd4}: kernel_rom_out = 16'sd16781;
            {4'd7, 3'd7, 3'd5}: kernel_rom_out = -16'sd7665;
            {4'd7, 3'd7, 3'd6}: kernel_rom_out = -16'sd122;
            {4'd7, 3'd7, 3'd7}: kernel_rom_out = 16'sd1083;

            // MODE 8: RFT-MANIFOLD (unitarity: 2.26e-15)
            {4'd8, 3'd0, 3'd0}: kernel_rom_out = -16'sd9374;
            {4'd8, 3'd0, 3'd1}: kernel_rom_out = -16'sd14997;
            {4'd8, 3'd0, 3'd2}: kernel_rom_out = -16'sd10409;
            {4'd8, 3'd0, 3'd3}: kernel_rom_out = -16'sd14601;
            {4'd8, 3'd0, 3'd4}: kernel_rom_out = -16'sd2148;
            {4'd8, 3'd0, 3'd5}: kernel_rom_out = -16'sd6335;
            {4'd8, 3'd0, 3'd6}: kernel_rom_out = -16'sd7654;
            {4'd8, 3'd0, 3'd7}: kernel_rom_out = 16'sd18330;
            {4'd8, 3'd1, 3'd0}: kernel_rom_out = -16'sd15451;
            {4'd8, 3'd1, 3'd1}: kernel_rom_out = -16'sd2699;
            {4'd8, 3'd1, 3'd2}: kernel_rom_out = 16'sd14530;
            {4'd8, 3'd1, 3'd3}: kernel_rom_out = -16'sd4158;
            {4'd8, 3'd1, 3'd4}: kernel_rom_out = 16'sd9216;
            {4'd8, 3'd1, 3'd5}: kernel_rom_out = -16'sd9076;
            {4'd8, 3'd1, 3'd6}: kernel_rom_out = 16'sd20734;
            {4'd8, 3'd1, 3'd7}: kernel_rom_out = 16'sd1429;
            {4'd8, 3'd2, 3'd0}: kernel_rom_out = -16'sd13688;
            {4'd8, 3'd2, 3'd1}: kernel_rom_out = 16'sd9764;
            {4'd8, 3'd2, 3'd2}: kernel_rom_out = -16'sd12176;
            {4'd8, 3'd2, 3'd3}: kernel_rom_out = 16'sd2159;
            {4'd8, 3'd2, 3'd4}: kernel_rom_out = -16'sd1565;
            {4'd8, 3'd2, 3'd5}: kernel_rom_out = -16'sd19719;
            {4'd8, 3'd2, 3'd6}: kernel_rom_out = -16'sd6927;
            {4'd8, 3'd2, 3'd7}: kernel_rom_out = -16'sd14099;
            {4'd8, 3'd3, 3'd0}: kernel_rom_out = -16'sd4780;
            {4'd8, 3'd3, 3'd1}: kernel_rom_out = 16'sd14468;
            {4'd8, 3'd3, 3'd2}: kernel_rom_out = 16'sd8313;
            {4'd8, 3'd3, 3'd3}: kernel_rom_out = -16'sd17369;
            {4'd8, 3'd3, 3'd4}: kernel_rom_out = -16'sd21091;
            {4'd8, 3'd3, 3'd5}: kernel_rom_out = 16'sd5047;
            {4'd8, 3'd3, 3'd6}: kernel_rom_out = 16'sd609;
            {4'd8, 3'd3, 3'd7}: kernel_rom_out = -16'sd196;
            {4'd8, 3'd4, 3'd0}: kernel_rom_out = 16'sd4780;
            {4'd8, 3'd4, 3'd1}: kernel_rom_out = 16'sd14468;
            {4'd8, 3'd4, 3'd2}: kernel_rom_out = -16'sd8313;
            {4'd8, 3'd4, 3'd3}: kernel_rom_out = -16'sd17369;
            {4'd8, 3'd4, 3'd4}: kernel_rom_out = 16'sd21091;
            {4'd8, 3'd4, 3'd5}: kernel_rom_out = 16'sd5047;
            {4'd8, 3'd4, 3'd6}: kernel_rom_out = 16'sd609;
            {4'd8, 3'd4, 3'd7}: kernel_rom_out = 16'sd196;
            {4'd8, 3'd5, 3'd0}: kernel_rom_out = 16'sd13688;
            {4'd8, 3'd5, 3'd1}: kernel_rom_out = 16'sd9764;
            {4'd8, 3'd5, 3'd2}: kernel_rom_out = 16'sd12176;
            {4'd8, 3'd5, 3'd3}: kernel_rom_out = 16'sd2159;
            {4'd8, 3'd5, 3'd4}: kernel_rom_out = 16'sd1565;
            {4'd8, 3'd5, 3'd5}: kernel_rom_out = -16'sd19719;
            {4'd8, 3'd5, 3'd6}: kernel_rom_out = -16'sd6927;
            {4'd8, 3'd5, 3'd7}: kernel_rom_out = 16'sd14099;
            {4'd8, 3'd6, 3'd0}: kernel_rom_out = 16'sd15451;
            {4'd8, 3'd6, 3'd1}: kernel_rom_out = -16'sd2699;
            {4'd8, 3'd6, 3'd2}: kernel_rom_out = -16'sd14530;
            {4'd8, 3'd6, 3'd3}: kernel_rom_out = -16'sd4158;
            {4'd8, 3'd6, 3'd4}: kernel_rom_out = -16'sd9216;
            {4'd8, 3'd6, 3'd5}: kernel_rom_out = -16'sd9076;
            {4'd8, 3'd6, 3'd6}: kernel_rom_out = 16'sd20734;
            {4'd8, 3'd6, 3'd7}: kernel_rom_out = -16'sd1429;
            {4'd8, 3'd7, 3'd0}: kernel_rom_out = 16'sd9374;
            {4'd8, 3'd7, 3'd1}: kernel_rom_out = -16'sd14997;
            {4'd8, 3'd7, 3'd2}: kernel_rom_out = 16'sd10409;
            {4'd8, 3'd7, 3'd3}: kernel_rom_out = -16'sd14601;
            {4'd8, 3'd7, 3'd4}: kernel_rom_out = 16'sd2148;
            {4'd8, 3'd7, 3'd5}: kernel_rom_out = -16'sd6335;
            {4'd8, 3'd7, 3'd6}: kernel_rom_out = -16'sd7654;
            {4'd8, 3'd7, 3'd7}: kernel_rom_out = -16'sd18330;

            // MODE 9: RFT-EULER (unitarity: 3.02e-15)
            {4'd9, 3'd0, 3'd0}: kernel_rom_out = -16'sd16232;
            {4'd9, 3'd0, 3'd1}: kernel_rom_out = 16'sd5203;
            {4'd9, 3'd0, 3'd2}: kernel_rom_out = -16'sd3776;
            {4'd9, 3'd0, 3'd3}: kernel_rom_out = -16'sd11809;
            {4'd9, 3'd0, 3'd4}: kernel_rom_out = 16'sd19982;
            {4'd9, 3'd0, 3'd5}: kernel_rom_out = -16'sd4049;
            {4'd9, 3'd0, 3'd6}: kernel_rom_out = 16'sd9809;
            {4'd9, 3'd0, 3'd7}: kernel_rom_out = -16'sd10839;
            {4'd9, 3'd1, 3'd0}: kernel_rom_out = -16'sd2338;
            {4'd9, 3'd1, 3'd1}: kernel_rom_out = 16'sd18201;
            {4'd9, 3'd1, 3'd2}: kernel_rom_out = -16'sd5501;
            {4'd9, 3'd1, 3'd3}: kernel_rom_out = -16'sd14165;
            {4'd9, 3'd1, 3'd4}: kernel_rom_out = -16'sd10024;
            {4'd9, 3'd1, 3'd5}: kernel_rom_out = 16'sd9963;
            {4'd9, 3'd1, 3'd6}: kernel_rom_out = 16'sd8648;
            {4'd9, 3'd1, 3'd7}: kernel_rom_out = 16'sd15213;
            {4'd9, 3'd2, 3'd0}: kernel_rom_out = 16'sd13633;
            {4'd9, 3'd2, 3'd1}: kernel_rom_out = 16'sd7122;
            {4'd9, 3'd2, 3'd2}: kernel_rom_out = -16'sd12391;
            {4'd9, 3'd2, 3'd3}: kernel_rom_out = -16'sd13010;
            {4'd9, 3'd2, 3'd4}: kernel_rom_out = 16'sd4481;
            {4'd9, 3'd2, 3'd5}: kernel_rom_out = -16'sd13424;
            {4'd9, 3'd2, 3'd6}: kernel_rom_out = -16'sd17677;
            {4'd9, 3'd2, 3'd7}: kernel_rom_out = -16'sd1227;
            {4'd9, 3'd3, 3'd0}: kernel_rom_out = 16'sd9056;
            {4'd9, 3'd3, 3'd1}: kernel_rom_out = -16'sd11303;
            {4'd9, 3'd3, 3'd2}: kernel_rom_out = -16'sd18406;
            {4'd9, 3'd3, 3'd3}: kernel_rom_out = -16'sd5239;
            {4'd9, 3'd3, 3'd4}: kernel_rom_out = -16'sd4120;
            {4'd9, 3'd3, 3'd5}: kernel_rom_out = 16'sd15523;
            {4'd9, 3'd3, 3'd6}: kernel_rom_out = 16'sd7303;
            {4'd9, 3'd3, 3'd7}: kernel_rom_out = -16'sd13653;
            {4'd9, 3'd4, 3'd0}: kernel_rom_out = -16'sd9056;
            {4'd9, 3'd4, 3'd1}: kernel_rom_out = -16'sd11303;
            {4'd9, 3'd4, 3'd2}: kernel_rom_out = -16'sd18406;
            {4'd9, 3'd4, 3'd3}: kernel_rom_out = 16'sd5239;
            {4'd9, 3'd4, 3'd4}: kernel_rom_out = -16'sd4120;
            {4'd9, 3'd4, 3'd5}: kernel_rom_out = -16'sd15523;
            {4'd9, 3'd4, 3'd6}: kernel_rom_out = 16'sd7303;
            {4'd9, 3'd4, 3'd7}: kernel_rom_out = 16'sd13653;
            {4'd9, 3'd5, 3'd0}: kernel_rom_out = -16'sd13633;
            {4'd9, 3'd5, 3'd1}: kernel_rom_out = 16'sd7122;
            {4'd9, 3'd5, 3'd2}: kernel_rom_out = -16'sd12391;
            {4'd9, 3'd5, 3'd3}: kernel_rom_out = 16'sd13010;
            {4'd9, 3'd5, 3'd4}: kernel_rom_out = 16'sd4481;
            {4'd9, 3'd5, 3'd5}: kernel_rom_out = 16'sd13424;
            {4'd9, 3'd5, 3'd6}: kernel_rom_out = -16'sd17677;
            {4'd9, 3'd5, 3'd7}: kernel_rom_out = 16'sd1227;
            {4'd9, 3'd6, 3'd0}: kernel_rom_out = 16'sd2338;
            {4'd9, 3'd6, 3'd1}: kernel_rom_out = 16'sd18201;
            {4'd9, 3'd6, 3'd2}: kernel_rom_out = -16'sd5501;
            {4'd9, 3'd6, 3'd3}: kernel_rom_out = 16'sd14165;
            {4'd9, 3'd6, 3'd4}: kernel_rom_out = -16'sd10024;
            {4'd9, 3'd6, 3'd5}: kernel_rom_out = -16'sd9963;
            {4'd9, 3'd6, 3'd6}: kernel_rom_out = 16'sd8648;
            {4'd9, 3'd6, 3'd7}: kernel_rom_out = -16'sd15213;
            {4'd9, 3'd7, 3'd0}: kernel_rom_out = 16'sd16232;
            {4'd9, 3'd7, 3'd1}: kernel_rom_out = 16'sd5203;
            {4'd9, 3'd7, 3'd2}: kernel_rom_out = -16'sd3776;
            {4'd9, 3'd7, 3'd3}: kernel_rom_out = 16'sd11809;
            {4'd9, 3'd7, 3'd4}: kernel_rom_out = 16'sd19982;
            {4'd9, 3'd7, 3'd5}: kernel_rom_out = 16'sd4049;
            {4'd9, 3'd7, 3'd6}: kernel_rom_out = 16'sd9809;
            {4'd9, 3'd7, 3'd7}: kernel_rom_out = 16'sd10839;

            // MODE 10: RFT-PHASE_COH (unitarity: 3.36e-15)
            {4'd10, 3'd0, 3'd0}: kernel_rom_out = -16'sd11229;
            {4'd10, 3'd0, 3'd1}: kernel_rom_out = -16'sd15554;
            {4'd10, 3'd0, 3'd2}: kernel_rom_out = 16'sd5617;
            {4'd10, 3'd0, 3'd3}: kernel_rom_out = -16'sd13614;
            {4'd10, 3'd0, 3'd4}: kernel_rom_out = -16'sd14765;
            {4'd10, 3'd0, 3'd5}: kernel_rom_out = 16'sd2171;
            {4'd10, 3'd0, 3'd6}: kernel_rom_out = 16'sd10240;
            {4'd10, 3'd0, 3'd7}: kernel_rom_out = 16'sd12696;
            {4'd10, 3'd1, 3'd0}: kernel_rom_out = -16'sd11768;
            {4'd10, 3'd1, 3'd1}: kernel_rom_out = 16'sd6617;
            {4'd10, 3'd1, 3'd2}: kernel_rom_out = -16'sd14607;
            {4'd10, 3'd1, 3'd3}: kernel_rom_out = -16'sd16824;
            {4'd10, 3'd1, 3'd4}: kernel_rom_out = 16'sd10658;
            {4'd10, 3'd1, 3'd5}: kernel_rom_out = 16'sd5380;
            {4'd10, 3'd1, 3'd6}: kernel_rom_out = -16'sd13456;
            {4'd10, 3'd1, 3'd7}: kernel_rom_out = 16'sd8449;
            {4'd10, 3'd2, 3'd0}: kernel_rom_out = -16'sd11428;
            {4'd10, 3'd2, 3'd1}: kernel_rom_out = 16'sd5462;
            {4'd10, 3'd2, 3'd2}: kernel_rom_out = 16'sd15937;
            {4'd10, 3'd2, 3'd3}: kernel_rom_out = -16'sd7178;
            {4'd10, 3'd2, 3'd4}: kernel_rom_out = 16'sd11876;
            {4'd10, 3'd2, 3'd5}: kernel_rom_out = -16'sd21097;
            {4'd10, 3'd2, 3'd6}: kernel_rom_out = 16'sd3226;
            {4'd10, 3'd2, 3'd7}: kernel_rom_out = -16'sd3346;
            {4'd10, 3'd3, 3'd0}: kernel_rom_out = -16'sd11902;
            {4'd10, 3'd3, 3'd1}: kernel_rom_out = -16'sd14876;
            {4'd10, 3'd3, 3'd2}: kernel_rom_out = -16'sd6159;
            {4'd10, 3'd3, 3'd3}: kernel_rom_out = 16'sd4114;
            {4'd10, 3'd3, 3'd4}: kernel_rom_out = -16'sd8012;
            {4'd10, 3'd3, 3'd5}: kernel_rom_out = -16'sd7623;
            {4'd10, 3'd3, 3'd6}: kernel_rom_out = -16'sd15508;
            {4'd10, 3'd3, 3'd7}: kernel_rom_out = -16'sd17119;
            {4'd10, 3'd4, 3'd0}: kernel_rom_out = -16'sd11902;
            {4'd10, 3'd4, 3'd1}: kernel_rom_out = 16'sd14876;
            {4'd10, 3'd4, 3'd2}: kernel_rom_out = -16'sd6159;
            {4'd10, 3'd4, 3'd3}: kernel_rom_out = -16'sd4114;
            {4'd10, 3'd4, 3'd4}: kernel_rom_out = -16'sd8012;
            {4'd10, 3'd4, 3'd5}: kernel_rom_out = 16'sd7623;
            {4'd10, 3'd4, 3'd6}: kernel_rom_out = 16'sd15508;
            {4'd10, 3'd4, 3'd7}: kernel_rom_out = -16'sd17119;
            {4'd10, 3'd5, 3'd0}: kernel_rom_out = -16'sd11428;
            {4'd10, 3'd5, 3'd1}: kernel_rom_out = -16'sd5462;
            {4'd10, 3'd5, 3'd2}: kernel_rom_out = 16'sd15937;
            {4'd10, 3'd5, 3'd3}: kernel_rom_out = 16'sd7178;
            {4'd10, 3'd5, 3'd4}: kernel_rom_out = 16'sd11876;
            {4'd10, 3'd5, 3'd5}: kernel_rom_out = 16'sd21097;
            {4'd10, 3'd5, 3'd6}: kernel_rom_out = -16'sd3226;
            {4'd10, 3'd5, 3'd7}: kernel_rom_out = -16'sd3346;
            {4'd10, 3'd6, 3'd0}: kernel_rom_out = -16'sd11768;
            {4'd10, 3'd6, 3'd1}: kernel_rom_out = -16'sd6617;
            {4'd10, 3'd6, 3'd2}: kernel_rom_out = -16'sd14607;
            {4'd10, 3'd6, 3'd3}: kernel_rom_out = 16'sd16824;
            {4'd10, 3'd6, 3'd4}: kernel_rom_out = 16'sd10658;
            {4'd10, 3'd6, 3'd5}: kernel_rom_out = -16'sd5380;
            {4'd10, 3'd6, 3'd6}: kernel_rom_out = 16'sd13456;
            {4'd10, 3'd6, 3'd7}: kernel_rom_out = 16'sd8449;
            {4'd10, 3'd7, 3'd0}: kernel_rom_out = -16'sd11229;
            {4'd10, 3'd7, 3'd1}: kernel_rom_out = 16'sd15554;
            {4'd10, 3'd7, 3'd2}: kernel_rom_out = 16'sd5617;
            {4'd10, 3'd7, 3'd3}: kernel_rom_out = 16'sd13614;
            {4'd10, 3'd7, 3'd4}: kernel_rom_out = -16'sd14765;
            {4'd10, 3'd7, 3'd5}: kernel_rom_out = -16'sd2171;
            {4'd10, 3'd7, 3'd6}: kernel_rom_out = -16'sd10240;
            {4'd10, 3'd7, 3'd7}: kernel_rom_out = 16'sd12696;

            // MODE 11: RFT-ENTROPY (unitarity: 1.80e-15)
            {4'd11, 3'd0, 3'd0}: kernel_rom_out = -16'sd14051;
            {4'd11, 3'd0, 3'd1}: kernel_rom_out = -16'sd2494;
            {4'd11, 3'd0, 3'd2}: kernel_rom_out = 16'sd18787;
            {4'd11, 3'd0, 3'd3}: kernel_rom_out = -16'sd9991;
            {4'd11, 3'd0, 3'd4}: kernel_rom_out = -16'sd4227;
            {4'd11, 3'd0, 3'd5}: kernel_rom_out = -16'sd14890;
            {4'd11, 3'd0, 3'd6}: kernel_rom_out = 16'sd11475;
            {4'd11, 3'd0, 3'd7}: kernel_rom_out = -16'sd6781;
            {4'd11, 3'd1, 3'd0}: kernel_rom_out = -16'sd1723;
            {4'd11, 3'd1, 3'd1}: kernel_rom_out = -16'sd16243;
            {4'd11, 3'd1, 3'd2}: kernel_rom_out = 16'sd4200;
            {4'd11, 3'd1, 3'd3}: kernel_rom_out = 16'sd20030;
            {4'd11, 3'd1, 3'd4}: kernel_rom_out = -16'sd1295;
            {4'd11, 3'd1, 3'd5}: kernel_rom_out = -16'sd11445;
            {4'd11, 3'd1, 3'd6}: kernel_rom_out = -16'sd14446;
            {4'd11, 3'd1, 3'd7}: kernel_rom_out = -16'sd6833;
            {4'd11, 3'd2, 3'd0}: kernel_rom_out = 16'sd14915;
            {4'd11, 3'd2, 3'd1}: kernel_rom_out = -16'sd6872;
            {4'd11, 3'd2, 3'd2}: kernel_rom_out = -16'sd12760;
            {4'd11, 3'd2, 3'd3}: kernel_rom_out = -16'sd3770;
            {4'd11, 3'd2, 3'd4}: kernel_rom_out = -16'sd15825;
            {4'd11, 3'd2, 3'd5}: kernel_rom_out = -16'sd7052;
            {4'd11, 3'd2, 3'd6}: kernel_rom_out = 16'sd10854;
            {4'd11, 3'd2, 3'd7}: kernel_rom_out = -16'sd14456;
            {4'd11, 3'd3, 3'd0}: kernel_rom_out = 16'sd10675;
            {4'd11, 3'd3, 3'd1}: kernel_rom_out = 16'sd14818;
            {4'd11, 3'd3, 3'd2}: kernel_rom_out = 16'sd1849;
            {4'd11, 3'd3, 3'd3}: kernel_rom_out = -16'sd4649;
            {4'd11, 3'd3, 3'd4}: kernel_rom_out = 16'sd16336;
            {4'd11, 3'd3, 3'd5}: kernel_rom_out = -16'sd11593;
            {4'd11, 3'd3, 3'd6}: kernel_rom_out = -16'sd8869;
            {4'd11, 3'd3, 3'd7}: kernel_rom_out = -16'sd15336;
            {4'd11, 3'd4, 3'd0}: kernel_rom_out = -16'sd10675;
            {4'd11, 3'd4, 3'd1}: kernel_rom_out = 16'sd14818;
            {4'd11, 3'd4, 3'd2}: kernel_rom_out = 16'sd1849;
            {4'd11, 3'd4, 3'd3}: kernel_rom_out = 16'sd4649;
            {4'd11, 3'd4, 3'd4}: kernel_rom_out = -16'sd16336;
            {4'd11, 3'd4, 3'd5}: kernel_rom_out = 16'sd11593;
            {4'd11, 3'd4, 3'd6}: kernel_rom_out = -16'sd8869;
            {4'd11, 3'd4, 3'd7}: kernel_rom_out = -16'sd15336;
            {4'd11, 3'd5, 3'd0}: kernel_rom_out = -16'sd14915;
            {4'd11, 3'd5, 3'd1}: kernel_rom_out = -16'sd6872;
            {4'd11, 3'd5, 3'd2}: kernel_rom_out = -16'sd12760;
            {4'd11, 3'd5, 3'd3}: kernel_rom_out = 16'sd3770;
            {4'd11, 3'd5, 3'd4}: kernel_rom_out = 16'sd15825;
            {4'd11, 3'd5, 3'd5}: kernel_rom_out = 16'sd7052;
            {4'd11, 3'd5, 3'd6}: kernel_rom_out = 16'sd10854;
            {4'd11, 3'd5, 3'd7}: kernel_rom_out = -16'sd14456;
            {4'd11, 3'd6, 3'd0}: kernel_rom_out = 16'sd1723;
            {4'd11, 3'd6, 3'd1}: kernel_rom_out = -16'sd16243;
            {4'd11, 3'd6, 3'd2}: kernel_rom_out = 16'sd4200;
            {4'd11, 3'd6, 3'd3}: kernel_rom_out = -16'sd20030;
            {4'd11, 3'd6, 3'd4}: kernel_rom_out = 16'sd1295;
            {4'd11, 3'd6, 3'd5}: kernel_rom_out = 16'sd11445;
            {4'd11, 3'd6, 3'd6}: kernel_rom_out = -16'sd14446;
            {4'd11, 3'd6, 3'd7}: kernel_rom_out = -16'sd6833;
            {4'd11, 3'd7, 3'd0}: kernel_rom_out = 16'sd14051;
            {4'd11, 3'd7, 3'd1}: kernel_rom_out = -16'sd2494;
            {4'd11, 3'd7, 3'd2}: kernel_rom_out = 16'sd18787;
            {4'd11, 3'd7, 3'd3}: kernel_rom_out = 16'sd9991;
            {4'd11, 3'd7, 3'd4}: kernel_rom_out = 16'sd4227;
            {4'd11, 3'd7, 3'd5}: kernel_rom_out = 16'sd14890;
            {4'd11, 3'd7, 3'd6}: kernel_rom_out = 16'sd11475;
            {4'd11, 3'd7, 3'd7}: kernel_rom_out = -16'sd6781;
