// ===============================================
// QUANTONIUMOS FULL ENGINES - INTEGRATED DESIGN
// Combines RFT + Feistel-48 + SIS Hash + Compression Engines
// Based on canonical_true_rft.py, rft_sis_hash_v31.py, and feistel_48.c
// ===============================================
// SPDX-License-Identifier: LicenseRef-QuantoniumOS-Claims-NC
// Copyright (C) 2025 Luis M. Minier
// NOTE: Use .sv extension for SystemVerilog synthesis

`timescale 1ns/1ps
`default_nettype none  // Catch typos and undefined signals

// ===============================================
// ENGINE 1: CANONICAL RFT CORE
// Implements unitary RFT with golden-ratio parameterization
// Ψ = Σ_i w_i D_φi C_σi D†_φi
// ===============================================
module canonical_rft_core #(
    parameter N = 64,               // Transform size
    parameter PRECISION = 32        // Fixed-point precision (Q16.16)
) (
    input wire clk,
    input wire reset,
    input wire start,
    input wire [N*PRECISION-1:0] signal_in,  // Packed: concatenated input signal
    output reg [N*PRECISION-1:0] signal_out, // Packed: concatenated RFT coefficients
    output reg valid,
    output reg done
);

    // Golden ratio φ = (1 + √5) / 2 ≈ 1.618034 in Q16.16
    localparam [PRECISION-1:0] PHI = 32'h0001_9E37;  // 1.618034 in Q16.16
    
    // Transform states
    localparam IDLE = 3'd0;
    localparam SETUP_CORDIC = 3'd1;
    localparam WAIT_CORDIC = 3'd2;
    localparam APPLY_KERNEL = 3'd3;
    localparam ORTHONORMALIZE = 3'd4;
    localparam OUTPUT = 3'd5;
    
    reg [2:0] state;
    integer row_idx, col_idx;
    
    // Precomputed golden-ratio phase sequence: φ_k = frac(k/φ)
    reg [PRECISION-1:0] phi_sequence [0:N-1];
    
    // RFT basis matrix (complex, stored as real/imag pairs)
    reg [PRECISION-1:0] rft_matrix_real [0:N-1][0:N-1];
    reg [PRECISION-1:0] rft_matrix_imag [0:N-1][0:N-1];
    
    // Unpacked internal signal arrays
    reg [PRECISION-1:0] signal_in_unpacked [0:N-1];
    reg [PRECISION-1:0] signal_out_unpacked [0:N-1];
    
    // CORDIC outputs for sin/cos
    wire [PRECISION-1:0] cordic_sin, cordic_cos;
    wire cordic_valid;
    reg cordic_start;
    reg [PRECISION-1:0] cordic_angle;
    
    // Internal computation registers
    reg [PRECISION-1:0] kernel_weight;
    reg [PRECISION-1:0] phase_term;
    reg [63:0] accumulator_real, accumulator_imag;
    
    // Initialize golden-ratio phase sequence
    integer i;
    initial begin
        for (i = 0; i < N; i = i + 1) begin
            // φ_k = frac(k/φ) - compute fractional part
            // Simplified: use (k * 0x9E37) >> 16 & 0xFFFF for fractional part
            phi_sequence[i] = (i * PHI) & 32'h0000_FFFF;
        end
        // Debug
        $display("Phi Sequence[0]: %h", phi_sequence[0]);
        $display("Phi Sequence[1]: %h", phi_sequence[1]);
    end
    
    // Compute Gaussian kernel weight: exp(-0.5 * ((i-j)/(σ*N))^2)
    // Simplified for hardware: use lookup table or approximation
    function [PRECISION-1:0] gaussian_weight;
        input [7:0] i, j;
        reg signed [15:0] diff;
        begin
            diff = {8'b0, i} - {8'b0, j};
            // Approximation: w ≈ 1 - |diff|/N for small kernels
            if (diff < 0) diff = -diff;
            gaussian_weight = (32'h0001_0000) - (({16'b0, diff} << 16) / N);
        end
    endfunction
    
    // Unpack input signal
    integer unpack_idx;
    always @(*) begin
        for (unpack_idx = 0; unpack_idx < N; unpack_idx = unpack_idx + 1) begin
            signal_in_unpacked[unpack_idx] = signal_in[unpack_idx*PRECISION +: PRECISION];
        end
    end
    
    // Pack output signal
    integer pack_idx;
    always @(*) begin
        for (pack_idx = 0; pack_idx < N; pack_idx = pack_idx + 1) begin
            signal_out[pack_idx*PRECISION +: PRECISION] = signal_out_unpacked[pack_idx];
        end
    end
    
    // Main RFT computation FSM
    integer rst_i;
    integer debug_cnt = 0;
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            row_idx <= 0;
            col_idx <= 0;
            valid <= 0;
            done <= 0;
            cordic_start <= 0;
            accumulator_real <= 0;
            accumulator_imag <= 0;
            for (rst_i = 0; rst_i < N; rst_i = rst_i + 1) begin
                signal_out_unpacked[rst_i] <= 0;
            end
        end else begin
            debug_cnt <= debug_cnt + 1;
            // Debug print
            if (debug_cnt < 20 || state != IDLE) $display("RFT State: %d, Start: %b, Row: %d, Col: %d", state, start, row_idx, col_idx);
            
            case (state)
                IDLE: begin
                    if (start) begin
                        state <= SETUP_CORDIC;
                        row_idx <= 0;
                        col_idx <= 0;
                        valid <= 0;
                        done <= 0;
                    end
                end
                
                SETUP_CORDIC: begin
                    // Closed-Form Φ-RFT: Ψ_jk = (1/√N) * exp(i * 2π * (β{j/φ} + 0.5σj²/N - jk/N))
                    // j = row_idx, k = col_idx
                    
                    // Amplitude: 1/√N (For N=64, 1/8 = 0.125 = 0x2000)
                    kernel_weight <= 32'h0000_2000;
                    
                    // Phase Calculation: angle = 2π * ({j/φ} + 0.5j²/N - jk/N)
                    // 2π in Q16.16 = 0x6487E
                    // We compute terms directly in radians to avoid precision loss
                    
                    cordic_angle <= (
                        (phi_sequence[row_idx] * 32'h6487E) >>> 16
                    ) + (
                        ((row_idx * row_idx * 32'h6487E) / (2 * N))
                    ) - (
                        ((row_idx * col_idx * 32'h6487E) / N)
                    );
                    
                    cordic_start <= 1;
                    state <= WAIT_CORDIC;
                end

                WAIT_CORDIC: begin
                    cordic_start <= 0;
                    
                    // Wait for CORDIC
                    if (cordic_valid) begin
                        // Store kernel matrix element with proper complex exponential
                        // K[i,j] = w * (cos(θ) + j*sin(θ))
                        rft_matrix_real[row_idx][col_idx] <= (kernel_weight * cordic_cos) >>> 16;
                        rft_matrix_imag[row_idx][col_idx] <= (kernel_weight * cordic_sin) >>> 16;
                    
                        // Advance matrix construction
                        if (col_idx == N-1) begin
                            col_idx <= 0;
                            if (row_idx == N-1) begin
                                state <= APPLY_KERNEL;
                                row_idx <= 0;
                            end else begin
                                row_idx <= row_idx + 1;
                                state <= SETUP_CORDIC;
                            end
                        end else begin
                            col_idx <= col_idx + 1;
                            state <= SETUP_CORDIC;
                        end
                    end
                end
                
                APPLY_KERNEL: begin
                    // FIX B: Pipelined MAC - one multiply-accumulate per cycle
                    // Apply RFT: y = Ψ^H * x
                    // Compute dot product incrementally
                    
                    if (col_idx == 0) begin
                        // Initialize accumulator for new row
                        accumulator_real <= 0;
                        accumulator_imag <= 0;
                    end
                    
                    // Single MAC operation per cycle
                    // Complex multiply: (a + jb) * x = ax + j(bx)
                    accumulator_real <= accumulator_real + 
                        (rft_matrix_real[row_idx][col_idx] * signal_in_unpacked[col_idx]);
                    accumulator_imag <= accumulator_imag + 
                        (rft_matrix_imag[row_idx][col_idx] * signal_in_unpacked[col_idx]);
                    
                    // Advance through matrix
                    if (col_idx == N-1) begin
                        // Row complete - store result (magnitude)
                        signal_out_unpacked[row_idx] <= accumulator_real[47:16];  // Q16.16 result
                        col_idx <= 0;
                        
                        if (row_idx == N-1) begin
                            state <= OUTPUT;
                        end else begin
                            row_idx <= row_idx + 1;
                        end
                    end else begin
                        col_idx <= col_idx + 1;
                    end
                end
                
                OUTPUT: begin
                    valid <= 1;
                    done <= 1;
                    state <= IDLE;
                end
                default: state <= IDLE;
            endcase
        end
    end

endmodule

// ===============================================
// CORDIC IP CORE for sin/cos computation
// Computes cos(θ) and sin(θ) in Q16.16 fixed-point
// ===============================================
module cordic_sincos #(
    parameter WIDTH = 32
) (
    input wire clk,
    input wire reset,
    input wire start,
    input wire [WIDTH-1:0] angle,  // Input angle in Q16.16 (0 to 2π mapped to 0 to 2^16)
    output reg [WIDTH-1:0] cos_out, // cos(θ) in Q16.16
    output reg [WIDTH-1:0] sin_out, // sin(θ) in Q16.16
    output reg valid
);
    // CORDIC algorithm implementation
    // Using 16 iterations for Q16.16 precision
    localparam ITERATIONS = 16;
    localparam K = 32'h00009B74; // CORDIC gain factor ≈ 0.6073 in Q16.16
    
    reg [4:0] iteration;
    reg [WIDTH-1:0] x, y, z;
    reg computing;
    
    // CORDIC atan table (Q16.16 format)
    reg [WIDTH-1:0] atan_table [0:15];
    initial begin
        atan_table[0]  = 32'h0000C910; // atan(2^-0) = 45°
        atan_table[1]  = 32'h000076B2; // atan(2^-1) = 26.565°
        atan_table[2]  = 32'h00003EB7; // atan(2^-2)
        atan_table[3]  = 32'h00001FD6; // atan(2^-3)
        atan_table[4]  = 32'h00000FFB; // atan(2^-4)
        atan_table[5]  = 32'h000007FF; // atan(2^-5)
        atan_table[6]  = 32'h00000400; // atan(2^-6)
        atan_table[7]  = 32'h00000200; // atan(2^-7)
        atan_table[8]  = 32'h00000100; // atan(2^-8)
        atan_table[9]  = 32'h00000080; // atan(2^-9)
        atan_table[10] = 32'h00000040; // atan(2^-10)
        atan_table[11] = 32'h00000020; // atan(2^-11)
        atan_table[12] = 32'h00000010; // atan(2^-12)
        atan_table[13] = 32'h00000008; // atan(2^-13)
        atan_table[14] = 32'h00000004; // atan(2^-14)
        atan_table[15] = 32'h00000002; // atan(2^-15)
    end
    
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            computing <= 0;
            valid <= 0;
            iteration <= 0;
        end else if (start && !computing) begin
            // Initialize CORDIC
            x <= K; // Initial x = K (gain factor)
            y <= 0;
            z <= angle;
            iteration <= 0;
            computing <= 1;
            valid <= 0;
        end else if (computing) begin
            if (iteration < ITERATIONS) begin
                // CORDIC rotation
                if (z[WIDTH-1]) begin // z < 0
                    x <= x + (y >>> iteration);
                    y <= y - (x >>> iteration);
                    z <= z + atan_table[iteration];
                end else begin // z >= 0
                    x <= x - (y >>> iteration);
                    y <= y + (x >>> iteration);
                    z <= z - atan_table[iteration];
                end
                iteration <= iteration + 1;
            end else begin
                // Done
                cos_out <= x;
                sin_out <= y;
                valid <= 1;
                computing <= 0;
            end
        end else begin
            valid <= 0;
        end
    end
endmodule

// ===============================================
// ENGINE 2: RFT-SIS HASH v3.1 CORE
// Cryptographic coordinate expansion with SIS hardness
// ===============================================
module rft_sis_hash_v31 #(
    parameter SIS_N = 512,
    parameter SIS_M = 1024,
    parameter SIS_Q = 3329,
    parameter SIS_BETA = 100
) (
    input wire clk,
    input wire reset,
    input wire start,
    input wire [63:0] coordinate_x,     // Input coordinate (double precision bits)
    input wire [63:0] coordinate_y,
    input wire [63:0] coordinate_z,     // Optional 3D
    output reg [255:0] hash_digest,     // SHA3-256 output
    output reg valid
);

    // State machine
    localparam IDLE = 3'd0;
    localparam EXPAND_COORDS = 3'd1;
    localparam RFT_TRANSFORM = 3'd2;
    localparam SIS_QUANTIZE = 3'd3;
    localparam SIS_LATTICE = 3'd4;
    localparam HASH_FINAL = 3'd5;
    
    reg [2:0] state;
    integer loop_idx;
    
    // Expanded coordinate vector (cryptographic expansion)
    reg [63:0] expanded [0:SIS_N-1];
    
    // RFT output buffer
    reg [31:0] rft_output [0:SIS_N-1];
    
    // SIS quantized vector
    reg signed [15:0] sis_vector [0:SIS_N-1];
    
    // Lattice point accumulator
    reg signed [31:0] lattice_point [0:SIS_M-1];
    
    // SHA3 state (simplified interface - would need full SHA3 core)
    reg [1599:0] sha3_state;
    
    // Instantiate RFT core for coordinate transformation
    reg  [SIS_N*32-1:0] rft_signal_in_packed;
    wire [SIS_N*32-1:0] rft_signal_out_packed;
    wire rft_valid, rft_done;
    reg rft_start;
    
    // Pack/unpack helpers for RFT interface
    reg [31:0] rft_signal_in_array [0:SIS_N-1];
    reg [31:0] rft_signal_out_array [0:SIS_N-1];
    
    integer rft_pack_idx;
    always @(*) begin
        for (rft_pack_idx = 0; rft_pack_idx < SIS_N; rft_pack_idx = rft_pack_idx + 1) begin
            rft_signal_in_packed[rft_pack_idx*32 +: 32] = rft_signal_in_array[rft_pack_idx];
            rft_signal_out_array[rft_pack_idx] = rft_signal_out_packed[rft_pack_idx*32 +: 32];
        end
    end
    
    canonical_rft_core #(.N(SIS_N), .PRECISION(32)) rft_engine (
        .clk(clk),
        .reset(reset),
        .start(rft_start),
        .signal_in(rft_signal_in_packed),
        .signal_out(rft_signal_out_packed),
        .valid(rft_valid),
        .done(rft_done)
    );
    
    // FIX D: Cryptographic coordinate expansion
    // WARNING: Production requires SHAKE-128/256 XOF for secure sampling
    task expand_coordinates;
        input [63:0] x, y, z;
        integer i;
        reg [63:0] hash_state;
        begin
            // Stage 1: Direct coordinate embedding
            expanded[0] = x;
            expanded[1] = y;
            expanded[2] = z;
            
            // Stage 2: Cryptographic expansion (SIMPLIFIED - NOT SECURE)
            hash_state = x ^ y ^ z;
            for (i = 3; i < SIS_N; i = i + 1) begin
                // Davies-Meyer-like construction
                hash_state = hash_state ^ (expanded[i-1] + 64'h9E3779B97F4A7C15);
                hash_state = {hash_state[31:0], hash_state[63:32]} + hash_state; // Mix
                expanded[i] = hash_state;
            end
        end
    endtask
    
    // FIX D: SIS lattice matrix multiplication: As mod q
    // WARNING: Matrix A must be cryptographically generated in production
    task sis_lattice_multiply;
        integer i, j;
        reg signed [47:0] acc;
        reg [15:0] a_element;
        begin
            for (i = 0; i < SIS_M; i = i + 1) begin
                acc = 0;
                for (j = 0; j < SIS_N; j = j + 1) begin
                    // CRITICAL: Production needs SHAKE-128 generated matrix A
                    // Current: Deterministic placeholder (NOT secure)
                    a_element = 16'((i * 1103 + j * 3329 + 42) % SIS_Q);
                    acc = acc + (a_element * sis_vector[j]);
                end
                // Reduce mod q with proper signed handling
                lattice_point[i] = 32'(acc % SIS_Q);
                if (lattice_point[i] > (SIS_Q/2))
                    lattice_point[i] = lattice_point[i] - SIS_Q;
            end
        end
    endtask
    
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            valid <= 0;
            rft_start <= 0;
            hash_digest <= 0;
            for (loop_idx = 0; loop_idx < SIS_N; loop_idx = loop_idx + 1) begin
                expanded[loop_idx] <= 0;
                rft_output[loop_idx] <= 0;
                sis_vector[loop_idx] <= 0;
            end
            for (loop_idx = 0; loop_idx < SIS_M; loop_idx = loop_idx + 1) begin
                lattice_point[loop_idx] <= 0;
            end
        end else begin
            case (state)
                IDLE: begin
                    if (start) begin
                        state <= EXPAND_COORDS;
                        valid <= 0;
                    end
                end
                
                EXPAND_COORDS: begin
                    // FIX D: Cryptographically secure coordinate expansion
                    // WARNING: This is still simplified. Production needs SHAKE-128/256 XOF
                    expand_coordinates(coordinate_x, coordinate_y, coordinate_z);
                    
                    // Prepare RFT input
                    for (loop_idx = 0; loop_idx < SIS_N; loop_idx = loop_idx + 1) begin
                        rft_signal_in_array[loop_idx] = expanded[loop_idx][31:0];
                    end
                    
                    rft_start <= 1;
                    state <= RFT_TRANSFORM;
                end
                
                RFT_TRANSFORM: begin
                    rft_start <= 0;
                    if (rft_done) begin
                        // Capture RFT output
                        for (loop_idx = 0; loop_idx < SIS_N; loop_idx = loop_idx + 1) begin
                            rft_output[loop_idx] = rft_signal_out_array[loop_idx];
                        end
                        state <= SIS_QUANTIZE;
                    end
                end
                
                SIS_QUANTIZE: begin
                    // Quantize RFT output to SIS vector: s ∈ [-β, β]
                    for (loop_idx = 0; loop_idx < SIS_N; loop_idx = loop_idx + 1) begin
                        // Scale and clip to [-SIS_BETA, SIS_BETA]
                        sis_vector[loop_idx] = 16'(rft_output[loop_idx][30:16]) % SIS_BETA;
                    end
                    state <= SIS_LATTICE;
                end
                
                SIS_LATTICE: begin
                    // Compute lattice point: As mod q
                    sis_lattice_multiply();
                    state <= HASH_FINAL;
                end
                
                HASH_FINAL: begin
                    // FIX C: Real SHA3-256 (Keccak-f[1600]) needed here
                    // CRITICAL WARNING: This is NOT SHA3! 
                    // Production MUST use verified Keccak IP core from:
                    // - OpenCores Keccak (https://opencores.org/projects/sha3)
                    // - Xilinx Secure IP (for FPGA)
                    // - Cadence/Synopsys DesignWare (for ASIC)
                    //
                    // Current implementation is PLACEHOLDER ONLY:
                    hash_digest <= {lattice_point[7], lattice_point[6], 
                                   lattice_point[5], lattice_point[4],
                                   lattice_point[3], lattice_point[2],
                                   lattice_point[1], lattice_point[0]};
                    
                    // TODO: Replace above with:
                    // keccak_256 keccak (
                    //     .clk(clk), .reset(reset), .start(keccak_start),
                    //     .data_in(lattice_point_flattened),
                    //     .hash_out(hash_digest), .valid(keccak_valid)
                    // );
                    
                    valid <= 1;
                    state <= IDLE;
                end
                default: state <= IDLE;
            endcase
        end
    end

endmodule


// ===============================================
// ENGINE 3: FEISTEL-48 ROUND FUNCTION
// Based on feistel_48.c with AES S-box and MixColumns
// ===============================================
module feistel_round_function (
    input wire [63:0] right_in,         // 64-bit right half
    input wire [127:0] round_key,       // 128-bit round key
    output reg [63:0] f_output          // F-function output
);

    // AES S-box (first 64 entries for demo - full 256 in production)
    reg [7:0] SBOX [0:255];
    initial begin
        SBOX[  0] = 8'h63; SBOX[  1] = 8'h7C; SBOX[  2] = 8'h77; SBOX[  3] = 8'h7B;
        SBOX[  4] = 8'hF2; SBOX[  5] = 8'h6B; SBOX[  6] = 8'h6F; SBOX[  7] = 8'hC5;
        SBOX[  8] = 8'h30; SBOX[  9] = 8'h01; SBOX[ 10] = 8'h67; SBOX[ 11] = 8'h2B;
        SBOX[ 12] = 8'hFE; SBOX[ 13] = 8'hD7; SBOX[ 14] = 8'hAB; SBOX[ 15] = 8'h76;
        // ... (Full 256-entry S-box in production)
        SBOX[252] = 8'hB0; SBOX[253] = 8'h54; SBOX[254] = 8'hBB; SBOX[255] = 8'h16;
    end
    
    // Golden ratio constant φ for key mixing
    localparam [63:0] PHI_64 = 64'h9E3779B97F4A7C15;
    
    // F-function pipeline stages (now combinatorial)
    reg [63:0] stage1_xor;
    reg [63:0] stage2_sbox;
    reg [63:0] stage3_mix;
    reg [63:0] stage4_arx;
    
    always @(*) begin
        // Stage 1: XOR with round key
        stage1_xor = right_in ^ round_key[63:0];
        
        // Stage 2: Byte substitution (AES S-box)
        stage2_sbox[7:0]   = SBOX[stage1_xor[7:0]];
        stage2_sbox[15:8]  = SBOX[stage1_xor[15:8]];
        stage2_sbox[23:16] = SBOX[stage1_xor[23:16]];
        stage2_sbox[31:24] = SBOX[stage1_xor[31:24]];
        stage2_sbox[39:32] = SBOX[stage1_xor[39:32]];
        stage2_sbox[47:40] = SBOX[stage1_xor[47:40]];
        stage2_sbox[55:48] = SBOX[stage1_xor[55:48]];
        stage2_sbox[63:56] = SBOX[stage1_xor[63:56]];
        
        // Stage 3: MixColumns-style diffusion
        // Simplified: XOR with rotated copies
        stage3_mix = stage2_sbox ^ {stage2_sbox[6:0], stage2_sbox[63:7]} 
                                  ^ {stage2_sbox[10:0], stage2_sbox[63:11]};
        
        // Stage 4: ARX (Add-Rotate-XOR) with golden ratio
        stage4_arx = ((stage3_mix + PHI_64) ^ (stage3_mix <<< 13) ^ (stage3_mix >>> 29));
        
        // Final output
        f_output = stage4_arx ^ round_key[127:64];
        
        // Debug
        if (right_in != 0) $display("Feistel F: In=%h Key=%h Out=%h SBOX[0]=%h", right_in, round_key, f_output, SBOX[0]);
    end

endmodule


// ===============================================
// ENGINE 4: FEISTEL-48 CIPHER CONTROLLER
// 48 rounds with HKDF key schedule
// ===============================================
module feistel_48_cipher (
    input wire clk,
    input wire reset,
    input wire start,
    input wire encrypt_mode,            // 1=encrypt, 0=decrypt
    input wire [255:0] master_key,      // 256-bit master key
    input wire [127:0] plaintext,       // 128-bit block
    output reg [127:0] ciphertext,
    output reg done
);

    localparam ROUNDS = 48;
    // Deterministic constants for placeholder HKDF and whitening
    localparam [255:0] HKDF_SALT         = 256'h00112233445566778899AABBCCDDEEFF00112233445566778899AABBCCDDEEFF;
    localparam [255:0] PRE_WHITEN_CONST  = 256'hA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55A;
    localparam [255:0] POST_WHITEN_CONST = 256'h5AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA55AA5;
    
    // State machine
    localparam IDLE = 2'd0;
    localparam KEY_SCHEDULE = 2'd1;
    localparam PROCESSING = 2'd2;
    localparam DONE_STATE = 2'd3;
    
    reg [1:0] state;
    reg [5:0] round_counter;  // 0-47
    
    // Feistel state: 128-bit split into L/R
    reg [63:0] left, right;
    wire [63:0] f_out;
    reg [63:0] left_next, right_next;
    
    // Round keys (derived from master key)
    reg [127:0] round_keys [0:ROUNDS-1];
    reg [7:0] key_gen_idx;
    
    // Whitening keys
    reg [127:0] pre_whiten, post_whiten;
    
    // Instantiate F-function
    feistel_round_function f_func (
        .right_in(right),
        .round_key(round_keys[round_counter]),
        .f_output(f_out)
    );
    
    // FIX E: HKDF-based key derivation with HMAC-SHA256
    // WARNING: Production needs real HMAC-SHA256 IP core
    task derive_round_keys;
        input [255:0] mk;
        integer r;
        reg [255:0] prk;  // Pseudorandom key (HKDF extract)
        reg [127:0] okm;  // Output keying material (HKDF expand)
        reg [255:0] temp;
        begin
            // HKDF-Extract: PRK = HMAC-SHA256(salt, IKM)
            // Simplified: PRK = SHA256(salt || master_key)
            // Production MUST use real HMAC:
            prk = mk ^ HKDF_SALT;
            
            for (r = 0; r < ROUNDS; r = r + 1) begin
                // HKDF-Expand: OKM = HMAC-SHA256(PRK, info || counter)
                // Simplified: OKM = SHA256(PRK || info || r)
                // info = "RFT_ROUND_" || r || "_PHI"
                //
                // CRITICAL: Production needs verified HMAC-SHA256 IP:
                // - Xilinx HMAC IP core
                // - OpenCores sha256 + HMAC wrapper
                // - DesignWare Cryptographic IP
                //
                // Current placeholder:
                temp = prk ^ (r * 256'h9E3779B97F4A7C159E3779B97F4A7C15);
                temp = {temp[223:0], temp[255:224]} + temp;  // Mix
                okm = temp[127:0] ^ temp[255:128];
                round_keys[r] = okm;
            end
            
            // Derive whitening keys with domain separation
            temp = prk ^ PRE_WHITEN_CONST;
            pre_whiten = temp[127:0];
            temp = prk ^ POST_WHITEN_CONST;
            post_whiten = temp[255:128];
        end
    endtask
    
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            round_counter <= 0;
            done <= 0;
            ciphertext <= 0;
            left <= 0;
            right <= 0;
            left_next <= 0;
            right_next <= 0;
            pre_whiten <= 0;
            post_whiten <= 0;
            for (integer k=0; k<ROUNDS; k++) round_keys[k] <= 0;
        end else begin
            case (state)
                IDLE: begin
                    if (start) begin
                        state <= KEY_SCHEDULE;
                        key_gen_idx <= 0;
                        done <= 0;
                    end
                end
                
                KEY_SCHEDULE: begin
                    // Derive all round keys
                    derive_round_keys(master_key);
                    
                    // Initial whitening
                    left <= plaintext[127:64] ^ pre_whiten[127:64];
                    right <= plaintext[63:0] ^ pre_whiten[63:0];
                    
                    round_counter <= 0;
                    state <= PROCESSING;
                end
                
                PROCESSING: begin
                    // Feistel round: (L, R) -> (R, L ⊕ F(R, K))
                    left_next <= right;
                    right_next <= left ^ f_out;
                    
                    left <= left_next;
                    right <= right_next;
                    
                    if (round_counter == ROUNDS - 1) begin
                        // Final swap and whitening
                        ciphertext[127:64] <= right_next ^ post_whiten[127:64];
                        ciphertext[63:0] <= left_next ^ post_whiten[63:0];
                        state <= DONE_STATE;
                    end else begin
                        round_counter <= round_counter + 1;
                    end
                end
                
                DONE_STATE: begin
                    done <= 1;
                    state <= IDLE;
                end
                default: state <= IDLE;
            endcase
        end
    end

endmodule


// ===============================================
// ENGINE 5: UNIFIED QUANTONIUMOS CORE
// Integrates: RFT + RFT-SIS Hash + Feistel-48 + Compression
// ===============================================
module quantoniumos_unified_core #(
    parameter RFT_SIZE = 64,
    parameter SIS_N = 512,
    parameter FEISTEL_ROUNDS = 48
) (
    input wire clk,
    input wire reset,
    input wire start,
    input wire [2:0] mode,              // 0=RFT, 1=SIS_Hash, 2=Feistel, 3=Full_Pipeline
    input wire [255:0] master_key,
    input wire [127:0] data_in,
    output reg [255:0] data_out,        // Flexible output size
    output reg done,
    
    // Observability and metrics
    output wire [31:0] rft_energy,
    output wire [15:0] sis_collision_resistance,
    output wire [5:0] feistel_round_count,
    output wire [31:0] pipeline_throughput
);

    // Mode definitions
    localparam MODE_RFT_ONLY = 3'd0;
    localparam MODE_SIS_HASH = 3'd1;
    localparam MODE_FEISTEL = 3'd2;
    localparam MODE_FULL_PIPELINE = 3'd3;
    localparam MODE_COMPRESS = 3'd4;
    
    // Inter-engine signals (packed for module ports)
    reg [RFT_SIZE*32-1:0] rft_signal_in_packed;
    wire [RFT_SIZE*32-1:0] rft_signal_out_packed;
    reg [31:0] rft_signal_in_array [0:RFT_SIZE-1];
    reg [31:0] rft_signal_out_array [0:RFT_SIZE-1];
    wire rft_valid, rft_done;
    reg rft_start;
    
    // Pack/unpack RFT arrays
    integer rft_idx;
    always @(*) begin
        for (rft_idx = 0; rft_idx < RFT_SIZE; rft_idx = rft_idx + 1) begin
            rft_signal_in_packed[rft_idx*32 +: 32] = rft_signal_in_array[rft_idx];
            rft_signal_out_array[rft_idx] = rft_signal_out_packed[rft_idx*32 +: 32];
        end
    end
    
    wire [255:0] sis_hash_out;
    wire sis_hash_valid;
    reg sis_hash_start;
    
    wire [127:0] feistel_out;
    wire feistel_done;
    reg feistel_start;
    
    // Performance counters
    reg [31:0] cycle_counter;
    reg [31:0] throughput_accumulator;
    
    // Instantiate RFT Core
    canonical_rft_core #(
        .N(RFT_SIZE),
        .PRECISION(32)
    ) rft_engine (
        .clk(clk),
        .reset(reset),
        .start(rft_start),
        .signal_in(rft_signal_in_packed),
        .signal_out(rft_signal_out_packed),
        .valid(rft_valid),
        .done(rft_done)
    );
    
    // Instantiate RFT-SIS Hash
    rft_sis_hash_v31 #(
        .SIS_N(SIS_N),
        .SIS_M(1024),
        .SIS_Q(3329),
        .SIS_BETA(100)
    ) sis_hash_engine (
        .clk(clk),
        .reset(reset),
        .start(sis_hash_start),
        .coordinate_x(data_in[127:64]),
        .coordinate_y(data_in[63:0]),
        .coordinate_z(64'h0),
        .hash_digest(sis_hash_out),
        .valid(sis_hash_valid)
    );
    
    // Instantiate Feistel-48 Cipher
    feistel_48_cipher feistel_engine (
        .clk(clk),
        .reset(reset),
        .start(feistel_start),
        .encrypt_mode(1'b1),
        .master_key(master_key),
        .plaintext(data_in),
        .ciphertext(feistel_out),
        .done(feistel_done)
    );
    
    // Output observability
    assign rft_energy = rft_signal_out_array[0];  // Energy in first coefficient
    assign sis_collision_resistance = 16'hFFFF;  // Hardness indicator
    assign feistel_round_count = 6'd48;
    assign pipeline_throughput = throughput_accumulator;
    
    // Main control FSM
    reg [2:0] pipeline_stage;
    integer loop_i;
    
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            done <= 0;
            rft_start <= 0;
            sis_hash_start <= 0;
            feistel_start <= 0;
            cycle_counter <= 0;
            throughput_accumulator <= 0;
            pipeline_stage <= 0;
            data_out <= 256'h0;
            for (loop_i = 0; loop_i < RFT_SIZE; loop_i = loop_i + 1) begin
                rft_signal_in_array[loop_i] <= 0;
            end
        end else begin
            done <= 0;
            cycle_counter <= cycle_counter + 1;
            
            case (mode)
                MODE_RFT_ONLY: begin
                    // RFT transform only
                    if (start && !rft_start) begin
                        // Load input data into RFT signal
                        rft_signal_in_array[0] <= data_in[31:0];
                        rft_signal_in_array[1] <= data_in[63:32];
                        rft_signal_in_array[2] <= data_in[95:64];
                        rft_signal_in_array[3] <= data_in[127:96];
                        for (loop_i = 4; loop_i < RFT_SIZE; loop_i = loop_i + 1) begin
                            rft_signal_in_array[loop_i] <= 0;
                        end
                        rft_start <= 1;
                    end else begin
                        rft_start <= 0;
                    end
                    
                    if (rft_done) begin
                        data_out[31:0] <= rft_signal_out_array[0];
                        data_out[63:32] <= rft_signal_out_array[1];
                        data_out[95:64] <= rft_signal_out_array[2];
                        data_out[127:96] <= rft_signal_out_array[3];
                        done <= 1;
                        throughput_accumulator <= (128 * 1000000) / cycle_counter;
                    end
                end
                
                MODE_SIS_HASH: begin
                    // RFT-SIS hash only
                    if (start && !sis_hash_start) begin
                        sis_hash_start <= 1;
                    end else begin
                        sis_hash_start <= 0;
                    end
                    
                    if (sis_hash_valid) begin
                        data_out <= sis_hash_out;
                        done <= 1;
                        throughput_accumulator <= (256 * 1000000) / cycle_counter;
                    end
                end
                
                MODE_FEISTEL: begin
                    // Feistel-48 cipher only
                    if (start && !feistel_start) begin
                        feistel_start <= 1;
                    end else begin
                        feistel_start <= 0;
                    end
                    
                    if (feistel_done) begin
                        data_out[127:0] <= feistel_out;
                        done <= 1;
                        throughput_accumulator <= (128 * 1000000) / cycle_counter;
                    end
                end
                
                MODE_FULL_PIPELINE: begin
                    // Full pipeline: RFT → SIS Hash → Feistel → Output
                    case (pipeline_stage)
                        3'd0: begin
                            if (start) begin
                                rft_signal_in_array[0] <= data_in[31:0];
                                rft_signal_in_array[1] <= data_in[63:32];
                                rft_start <= 1;
                                pipeline_stage <= 3'd1;
                            end
                        end
                        
                        3'd1: begin
                            rft_start <= 0;
                            if (rft_done) begin
                                // Feed RFT output to SIS hash
                                sis_hash_start <= 1;
                                pipeline_stage <= 3'd2;
                            end
                        end
                        
                        3'd2: begin
                            sis_hash_start <= 0;
                            if (sis_hash_valid) begin
                                // Feed SIS hash to Feistel
                                feistel_start <= 1;
                                pipeline_stage <= 3'd3;
                            end
                        end
                        
                        3'd3: begin
                            feistel_start <= 0;
                            if (feistel_done) begin
                                data_out[127:0] <= feistel_out;
                                data_out[255:128] <= sis_hash_out[127:0];
                                done <= 1;
                                throughput_accumulator <= (256 * 1000000) / cycle_counter;
                                pipeline_stage <= 3'd0;
                            end
                        end
                        
                        default: pipeline_stage <= 3'd0;
                    endcase
                end
                
                default: begin
                    done <= 0;
                end
            endcase
        end
    end

endmodule
