// SPDX-License-Identifier: LicenseRef-QuantoniumOS-Claims-NC
// Copyright (C) 2025 Luis M. Minier / quantoniumos
//
// RFTPU Accelerator Testbench - Unit Tests for phi_rft_core
// ========================================================
// This testbench validates the RFT transform core against Python-generated
// golden vectors. It includes:
//   - Functional verification with known-good test vectors
//   - SVA properties for protocol and timing
//   - Coverage points for completeness
//   - Self-checking with tolerance-based comparison
//
// To run with Verilator:
//   verilator --binary -j 0 -Wall --trace \
//     -I../build -CFLAGS "-g" \
//     -top tb_rft_core tb_rft_core.sv ../build/rftpu_architecture.sv
//

`timescale 1ns/1ps

// Test vector include file (generated by rftpu_test_vectors.py)
`include "rft_test_vectors.svh"

module tb_rft_core;

  //=========================================================================
  // Parameters
  //=========================================================================
  localparam int CLK_PERIOD = 10;           // 100 MHz
  localparam int SAMPLE_WIDTH = 16;
  localparam int BLOCK_SAMPLES = 8;
  localparam int DIGEST_WIDTH = 256;
  localparam int CORE_LATENCY = 4;
  
  // Tolerance for fixed-point comparison (in LSBs)
  localparam int TOLERANCE = 128;  // ~0.4% tolerance for Q1.15

  //=========================================================================
  // Signals
  //=========================================================================
  logic clk = 0;
  logic rst_n;
  
  // RFT core interface
  logic [SAMPLE_WIDTH-1:0] sample_in [BLOCK_SAMPLES];
  logic                    start;
  logic [2:0]              mode;
  logic                    digest_valid;
  logic [DIGEST_WIDTH-1:0] digest_out;
  logic [15:0]             energy_out;
  logic                    cascade_mode;
  logic                    h3_enable;

  // Test tracking
  int test_count = 0;
  int pass_count = 0;
  int fail_count = 0;
  string current_test_name;

  //=========================================================================
  // Clock Generation
  //=========================================================================
  always #(CLK_PERIOD/2) clk = ~clk;

  //=========================================================================
  // DUT Instantiation - phi_rft_core
  //=========================================================================
  // Note: This requires the generated SystemVerilog from SandPiper
  // The phi_rft_core module is nested inside the TLV output
  
  // For standalone testing, we instantiate the core directly
  // In real integration, this would be part of rftpu_accelerator

  // Simplified interface wrapper (matches phi_rft_core ports)
  logic [127:0] sample_flat;
  logic [127:0] rft_real_out;
  logic [127:0] rft_imag_out;
  logic [15:0]  rft_real [BLOCK_SAMPLES];
  logic [15:0]  rft_imag [BLOCK_SAMPLES];

  // Pack samples into flat vector
  always_comb begin
    for (int i = 0; i < BLOCK_SAMPLES; i++) begin
      sample_flat[i*16 +: 16] = sample_in[i];
    end
  end
  
  // Unpack outputs
  always_comb begin
    for (int i = 0; i < BLOCK_SAMPLES; i++) begin
      rft_real[i] = rft_real_out[i*16 +: 16];
      rft_imag[i] = rft_imag_out[i*16 +: 16];
    end
  end

  // DUT: phi_rft_core (from rftpu_architecture.sv)
  // phi_rft_core #(
  //   .SAMPLE_WIDTH(SAMPLE_WIDTH),
  //   .BLOCK_SAMPLES(BLOCK_SAMPLES),
  //   .DIGEST_WIDTH(DIGEST_WIDTH)
  // ) dut (
  //   .clk(clk),
  //   .rst_n(rst_n),
  //   .sample_in(sample_flat),
  //   .start(start),
  //   .mode(mode),
  //   .digest_valid(digest_valid),
  //   .digest_out(digest_out),
  //   .energy_out(energy_out),
  //   .rft_real(rft_real_out),
  //   .rft_imag(rft_imag_out),
  //   .cascade_mode(cascade_mode),
  //   .h3_enable(h3_enable)
  // );

  // Behavioral model for standalone testing
  // (Replace with actual DUT when integrating)
  `ifdef USE_BEHAVIORAL_MODEL
    `include "rft_behavioral_model.svh"
  `else
    // Direct DUT connection goes here
  `endif

  //=========================================================================
  // Test Utilities
  //=========================================================================
  
  // Compare with tolerance
  function automatic bit compare_with_tolerance(
    input logic signed [15:0] actual,
    input logic signed [15:0] expected,
    input int tolerance
  );
    int diff;
    diff = $signed(actual) - $signed(expected);
    if (diff < 0) diff = -diff;
    return (diff <= tolerance);
  endfunction
  
  // Report test result
  task automatic report_test(
    input string name,
    input bit passed,
    input string details = ""
  );
    test_count++;
    if (passed) begin
      pass_count++;
      $display("[PASS] %s %s", name, details);
    end else begin
      fail_count++;
      $display("[FAIL] %s %s", name, details);
    end
  endtask
  
  // Wait for digest valid with timeout
  task automatic wait_digest_valid(input int timeout_cycles);
    int cycles = 0;
    while (!digest_valid && cycles < timeout_cycles) begin
      @(posedge clk);
      cycles++;
    end
    if (cycles >= timeout_cycles) begin
      $display("[ERROR] Timeout waiting for digest_valid");
    end
  endtask

  //=========================================================================
  // SVA Properties and Assertions
  //=========================================================================
  `ifndef VERILATOR  // Verilator has limited SVA support
  
  // Property: After start, digest_valid should appear within CORE_LATENCY+2 cycles
  property p_latency_bound;
    @(posedge clk) disable iff (!rst_n)
    start |-> ##[1:CORE_LATENCY+2] digest_valid;
  endproperty
  assert property (p_latency_bound) else
    $error("Latency exceeded: digest_valid not asserted within bound");
  
  // Property: digest_out should be stable when digest_valid is high
  property p_digest_stable;
    @(posedge clk) disable iff (!rst_n)
    digest_valid |-> ##1 (digest_valid && $stable(digest_out)) || !digest_valid;
  endproperty
  assert property (p_digest_stable) else
    $error("Digest not stable while valid");
  
  // Property: No start during active processing
  // (If we're still processing, another start is ignored)
  sequence s_processing;
    start ##[1:CORE_LATENCY] digest_valid;
  endsequence
  
  // Property: Energy output is non-negative (it's unsigned, so always true)
  property p_energy_valid;
    @(posedge clk) disable iff (!rst_n)
    digest_valid |-> (energy_out >= 0);
  endproperty
  assert property (p_energy_valid);
  
  `endif // VERILATOR

  //=========================================================================
  // Coverage Points
  //=========================================================================
  `ifndef VERILATOR
  
  covergroup cg_rft_modes @(posedge clk iff (start && rst_n));
    cp_mode: coverpoint mode {
      bins mode_0 = {0};
      bins mode_1 = {1};
      bins mode_2 = {2};
      bins mode_3 = {3};
      bins mode_others = {[4:7]};
    }
    
    cp_cascade: coverpoint cascade_mode {
      bins disabled = {0};
      bins enabled = {1};
    }
    
    cp_h3: coverpoint h3_enable {
      bins disabled = {0};
      bins enabled = {1};
    }
    
    // Cross coverage
    cx_mode_cascade: cross cp_mode, cp_cascade;
  endgroup
  
  covergroup cg_sample_values @(posedge clk iff (start && rst_n));
    // Cover interesting sample patterns
    cp_sample0: coverpoint sample_in[0][15:14] {
      bins zero = {2'b00};
      bins positive = {2'b01};
      bins negative = {2'b10, 2'b11};
    }
    
    // All-zero input
    cp_all_zero: coverpoint (sample_in[0] == 0 && sample_in[1] == 0 &&
                            sample_in[2] == 0 && sample_in[3] == 0 &&
                            sample_in[4] == 0 && sample_in[5] == 0 &&
                            sample_in[6] == 0 && sample_in[7] == 0) {
      bins all_zero = {1};
      bins not_all_zero = {0};
    }
  endgroup
  
  cg_rft_modes cov_modes;
  cg_sample_values cov_samples;
  
  initial begin
    cov_modes = new();
    cov_samples = new();
  end
  
  `endif // VERILATOR

  //=========================================================================
  // Test Stimulus
  //=========================================================================
  
  // Task: Run single RFT test vector
  task automatic run_rft_test(input int test_idx);
    bit test_passed;
    int diff;
    
    current_test_name = rft_test_names[test_idx];
    $display("\n--- Running RFT Test %0d: %s ---", test_idx, current_test_name);
    
    // Load input samples (real only for now, imag assumed 0)
    for (int i = 0; i < BLOCK_SAMPLES; i++) begin
      sample_in[i] = rft_test_input_real[test_idx][i];
    end
    
    // Configure mode
    mode = 3'b001;  // Standard RFT mode
    cascade_mode = 0;
    h3_enable = 0;
    
    // Apply start pulse
    @(posedge clk);
    start = 1;
    @(posedge clk);
    start = 0;
    
    // Wait for result
    wait_digest_valid(CORE_LATENCY + 10);
    
    // Check outputs
    test_passed = 1;
    for (int i = 0; i < BLOCK_SAMPLES; i++) begin
      // Compare real part
      if (!compare_with_tolerance(rft_real[i], rft_test_expected_real[test_idx][i], TOLERANCE)) begin
        diff = $signed(rft_real[i]) - $signed(rft_test_expected_real[test_idx][i]);
        $display("  Real[%0d] mismatch: got %h, expected %h (diff=%0d)", 
                 i, rft_real[i], rft_test_expected_real[test_idx][i], diff);
        test_passed = 0;
      end
      
      // Compare imag part
      if (!compare_with_tolerance(rft_imag[i], rft_test_expected_imag[test_idx][i], TOLERANCE)) begin
        diff = $signed(rft_imag[i]) - $signed(rft_test_expected_imag[test_idx][i]);
        $display("  Imag[%0d] mismatch: got %h, expected %h (diff=%0d)", 
                 i, rft_imag[i], rft_test_expected_imag[test_idx][i], diff);
        test_passed = 0;
      end
    end
    
    report_test(current_test_name, test_passed);
    
    // Small gap between tests
    repeat(2) @(posedge clk);
  endtask
  
  // Task: Run all RFT tests
  task automatic run_all_rft_tests();
    $display("\n========================================");
    $display("Running All RFT Test Vectors");
    $display("========================================");
    
    for (int i = 0; i < NUM_RFT_TESTS; i++) begin
      run_rft_test(i);
    end
  endtask
  
  // Task: Run edge case tests
  task automatic run_edge_case_tests();
    $display("\n========================================");
    $display("Running Edge Case Tests");
    $display("========================================");
    
    // Test: Back-to-back starts
    $display("\n--- Back-to-back start test ---");
    for (int i = 0; i < BLOCK_SAMPLES; i++) begin
      sample_in[i] = 16'h1000;
    end
    mode = 3'b001;
    
    @(posedge clk);
    start = 1;
    @(posedge clk);
    start = 0;
    wait_digest_valid(CORE_LATENCY + 5);
    
    // Immediately start next
    start = 1;
    @(posedge clk);
    start = 0;
    wait_digest_valid(CORE_LATENCY + 5);
    
    report_test("back_to_back", 1);  // Pass if no hang
    
    // Test: Reset during processing
    $display("\n--- Reset during processing ---");
    start = 1;
    @(posedge clk);
    start = 0;
    @(posedge clk);
    @(posedge clk);
    rst_n = 0;  // Assert reset mid-processing
    @(posedge clk);
    rst_n = 1;
    repeat(5) @(posedge clk);
    
    report_test("reset_recovery", !digest_valid);  // Should not be valid after reset
  endtask

  //=========================================================================
  // Main Test Sequence
  //=========================================================================
  initial begin
    $display("#######################################################");
    $display("# RFTPU Accelerator Testbench - RFT Core Validation #");
    $display("#######################################################");
    
    // Initialize
    rst_n = 0;
    start = 0;
    mode = 0;
    cascade_mode = 0;
    h3_enable = 0;
    for (int i = 0; i < BLOCK_SAMPLES; i++) begin
      sample_in[i] = 0;
    end
    
    // Reset sequence
    repeat(10) @(posedge clk);
    rst_n = 1;
    repeat(5) @(posedge clk);
    
    // Run test suites
    run_all_rft_tests();
    run_edge_case_tests();
    
    // Final report
    $display("\n######################################################");
    $display("# TEST SUMMARY                                       #");
    $display("######################################################");
    $display("  Total Tests: %0d", test_count);
    $display("  Passed:      %0d", pass_count);
    $display("  Failed:      %0d", fail_count);
    $display("######################################################\n");
    
    if (fail_count == 0) begin
      $display("*** ALL TESTS PASSED ***\n");
    end else begin
      $display("*** SOME TESTS FAILED ***\n");
    end
    
    // Coverage report
    `ifndef VERILATOR
    $display("Coverage: Modes=%0.1f%%, Samples=%0.1f%%",
             cov_modes.get_coverage(), cov_samples.get_coverage());
    `endif
    
    $finish;
  end

  //=========================================================================
  // Waveform Dump
  //=========================================================================
  initial begin
    `ifdef TRACE
    $dumpfile("tb_rft_core.vcd");
    $dumpvars(0, tb_rft_core);
    `endif
  end

endmodule
