// SPDX-License-Identifier: LicenseRef-QuantoniumOS-Claims-NC
// Copyright (C) 2025 Luis M. Minier / quantoniumos
// Patent Application: USPTO #19/169,399
//
// ═══════════════════════════════════════════════════════════════════════════
// QUANTONIUMOS RFTPU - ALL 12 PROVEN RFT TRANSFORMS
// ═══════════════════════════════════════════════════════════════════════════
// 
// This chip embodies the FULL computational stack of QuantoniumOS:
//
// OPERATOR-BASED TRANSFORMS (Eigenbasis of K = T(R·d)):
//   Mode 0: RFT-Golden      - Golden ratio resonance (PRIMARY)
//   Mode 1: RFT-Fibonacci   - Fibonacci frequency structure
//   Mode 2: RFT-Harmonic    - Natural harmonic overtones (audio/music)
//   Mode 3: RFT-Geometric   - Self-similar φ^i frequencies
//   Mode 4: RFT-Beating     - Golden ratio interference patterns
//   Mode 5: RFT-Phyllotaxis - Golden angle 137.5° (biological)
//   Mode 6: RFT-Cascade     - H3 DCT+RFT blend (universal compression)
//   Mode 7: RFT-Hybrid-DCT  - Split DCT/RFT basis (mixed content)
//
// PATENT VARIANTS (USPTO 19/169,399):
//   Mode 8:  RFT-Manifold   - Manifold projection (+47.9 dB winner)
//   Mode 9:  RFT-Euler      - Spherical geodesic resonance  
//   Mode 10: RFT-PhaseCoh   - Phase-space coherence (chirp signals)
//   Mode 11: RFT-Entropy    - Entropy-modulated chaos (noise-like)
//
// DEMO MODES:
//   Mode 12: SIS Hash       - Post-quantum lattice demo
//   Mode 13: Feistel-48     - Cipher demo
//   Mode 14: Quantum Sim    - GHZ state demo
//   Mode 15: Roundtrip      - Forward + inverse test
//
// All 12 RFT kernels: Q1.15 fixed-point, unitarity error < 1e-13
// Generated from: algorithms/rft/variants/operator_variants.py
// Cross-validated: Python reference matches RTL
//
// This file is listed in CLAIMS_PRACTICING_FILES.txt

/* verilator lint_off UNUSEDPARAM */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off WIDTHEXPAND */
/* verilator lint_off WIDTHTRUNC */

module fpga_top (
    input wire WF_CLK,
    input wire WF_BUTTON,
    output wire [7:0] WF_LED
);

    // Mode definitions
    localparam [3:0] MODE_RFT_GOLDEN      = 4'd0;
    localparam [3:0] MODE_RFT_FIBONACCI   = 4'd1;
    localparam [3:0] MODE_RFT_HARMONIC    = 4'd2;
    localparam [3:0] MODE_RFT_GEOMETRIC   = 4'd3;
    localparam [3:0] MODE_RFT_BEATING     = 4'd4;
    localparam [3:0] MODE_RFT_PHYLLOTAXIS = 4'd5;
    localparam [3:0] MODE_RFT_CASCADE     = 4'd6;
    localparam [3:0] MODE_RFT_HYBRID_DCT  = 4'd7;
    localparam [3:0] MODE_RFT_MANIFOLD    = 4'd8;
    localparam [3:0] MODE_RFT_EULER       = 4'd9;
    localparam [3:0] MODE_RFT_PHASE_COH   = 4'd10;
    localparam [3:0] MODE_RFT_ENTROPY     = 4'd11;
    localparam [3:0] MODE_SIS_HASH        = 4'd12;
    localparam [3:0] MODE_FEISTEL         = 4'd13;
    localparam [3:0] MODE_QUANTUM_SIM     = 4'd14;
    localparam [3:0] MODE_ROUNDTRIP       = 4'd15;

    // State machine
    localparam [2:0] STATE_IDLE    = 3'd0;
    localparam [2:0] STATE_COMPUTE = 3'd2;
    localparam [2:0] STATE_DONE    = 3'd5;

    // Registers
    reg [7:0] reset_counter = 8'h00;
    wire reset = (reset_counter < 8'd10);
    
    reg [19:0] button_debounce = 20'h00000;
    reg button_stable = 1'b0;
    reg button_prev = 1'b0;
    wire button_edge = button_stable && !button_prev;
    
    reg [3:0] current_mode = MODE_RFT_GOLDEN;
    reg [23:0] auto_cycle_counter = 24'h000000;
    wire auto_cycle_trigger = (auto_cycle_counter == 24'hFFFFFF);
    
    reg [7:0] cyc_cnt = 8'h00;
    wire start = button_edge || (cyc_cnt == 8'd20);
    
    reg [2:0] state = STATE_IDLE;
    reg [2:0] k_index = 3'b000;
    reg [2:0] n_index = 3'b000;
    
    reg [15:0] sample [0:7];
    reg valid = 1'b0;
    
    reg signed [15:0] kernel_reg;
    reg signed [15:0] kernel_rom_out;
    
    wire [15:0] input_selected = sample[n_index];
    wire signed [31:0] mult_out = $signed(input_selected) * $signed(kernel_reg);
    
    reg signed [31:0] acc = 32'sh00000000;
    reg signed [31:0] rft_out [0:7];
    
    wire is_computing = (state == STATE_COMPUTE);
    wire is_done = (state == STATE_DONE);
    wire save_result = (n_index == 3'b111) && is_computing;
    
    reg [7:0] led_output = 8'h00;
    
    integer i;

    // ═══════════════════════════════════════════════════════════════════════
    // KERNEL ROM: 12 kernels × 64 coefficients = 768 entries
    // ═══════════════════════════════════════════════════════════════════════
    
    always @(*) begin
        case ({current_mode, k_index, n_index})
// All 12 validated RFT kernels - case statement body
// Generated from algorithms/rft/variants/operator_variants.py

            // MODE 0: RFT-GOLDEN (unitarity: 6.12e-15)
            {4'd0, 3'd0, 3'd0}: kernel_rom_out = -16'sd10528;
            {4'd0, 3'd0, 3'd1}: kernel_rom_out = 16'sd12809;
            {4'd0, 3'd0, 3'd2}: kernel_rom_out = -16'sd11788;
            {4'd0, 3'd0, 3'd3}: kernel_rom_out = -16'sd12520;
            {4'd0, 3'd0, 3'd4}: kernel_rom_out = 16'sd14036;
            {4'd0, 3'd0, 3'd5}: kernel_rom_out = -16'sd14281;
            {4'd0, 3'd0, 3'd6}: kernel_rom_out = -16'sd9488;
            {4'd0, 3'd0, 3'd7}: kernel_rom_out = -16'sd3470;
            {4'd0, 3'd1, 3'd0}: kernel_rom_out = -16'sd11613;
            {4'd0, 3'd1, 3'd1}: kernel_rom_out = 16'sd12317;
            {4'd0, 3'd1, 3'd2}: kernel_rom_out = 16'sd11248;
            {4'd0, 3'd1, 3'd3}: kernel_rom_out = -16'sd7835;
            {4'd0, 3'd1, 3'd4}: kernel_rom_out = 16'sd9793;
            {4'd0, 3'd1, 3'd5}: kernel_rom_out = 16'sd15845;
            {4'd0, 3'd1, 3'd6}: kernel_rom_out = 16'sd13399;
            {4'd0, 3'd1, 3'd7}: kernel_rom_out = 16'sd8523;
            {4'd0, 3'd2, 3'd0}: kernel_rom_out = -16'sd12087;
            {4'd0, 3'd2, 3'd1}: kernel_rom_out = -16'sd10234;
            {4'd0, 3'd2, 3'd2}: kernel_rom_out = 16'sd11353;
            {4'd0, 3'd2, 3'd3}: kernel_rom_out = -16'sd15150;
            {4'd0, 3'd2, 3'd4}: kernel_rom_out = -16'sd8738;
            {4'd0, 3'd2, 3'd5}: kernel_rom_out = 16'sd7100;
            {4'd0, 3'd2, 3'd6}: kernel_rom_out = -16'sd13620;
            {4'd0, 3'd2, 3'd7}: kernel_rom_out = -16'sd12336;
            {4'd0, 3'd3, 3'd0}: kernel_rom_out = -16'sd12043;
            {4'd0, 3'd3, 3'd1}: kernel_rom_out = -16'sd10784;
            {4'd0, 3'd3, 3'd2}: kernel_rom_out = -16'sd11936;
            {4'd0, 3'd3, 3'd3}: kernel_rom_out = -16'sd9443;
            {4'd0, 3'd3, 3'd4}: kernel_rom_out = -16'sd12944;
            {4'd0, 3'd3, 3'd5}: kernel_rom_out = -16'sd5602;
            {4'd0, 3'd3, 3'd6}: kernel_rom_out = 16'sd9043;
            {4'd0, 3'd3, 3'd7}: kernel_rom_out = 16'sd17320;
            {4'd0, 3'd4, 3'd0}: kernel_rom_out = -16'sd12043;
            {4'd0, 3'd4, 3'd1}: kernel_rom_out = 16'sd10784;
            {4'd0, 3'd4, 3'd2}: kernel_rom_out = -16'sd11936;
            {4'd0, 3'd4, 3'd3}: kernel_rom_out = 16'sd9443;
            {4'd0, 3'd4, 3'd4}: kernel_rom_out = -16'sd12944;
            {4'd0, 3'd4, 3'd5}: kernel_rom_out = 16'sd5602;
            {4'd0, 3'd4, 3'd6}: kernel_rom_out = 16'sd9043;
            {4'd0, 3'd4, 3'd7}: kernel_rom_out = -16'sd17320;
            {4'd0, 3'd5, 3'd0}: kernel_rom_out = -16'sd12087;
            {4'd0, 3'd5, 3'd1}: kernel_rom_out = 16'sd10234;
            {4'd0, 3'd5, 3'd2}: kernel_rom_out = 16'sd11353;
            {4'd0, 3'd5, 3'd3}: kernel_rom_out = 16'sd15150;
            {4'd0, 3'd5, 3'd4}: kernel_rom_out = -16'sd8738;
            {4'd0, 3'd5, 3'd5}: kernel_rom_out = -16'sd7100;
            {4'd0, 3'd5, 3'd6}: kernel_rom_out = -16'sd13620;
            {4'd0, 3'd5, 3'd7}: kernel_rom_out = 16'sd12336;
            {4'd0, 3'd6, 3'd0}: kernel_rom_out = -16'sd11613;
            {4'd0, 3'd6, 3'd1}: kernel_rom_out = -16'sd12317;
            {4'd0, 3'd6, 3'd2}: kernel_rom_out = 16'sd11248;
            {4'd0, 3'd6, 3'd3}: kernel_rom_out = 16'sd7835;
            {4'd0, 3'd6, 3'd4}: kernel_rom_out = 16'sd9793;
            {4'd0, 3'd6, 3'd5}: kernel_rom_out = -16'sd15845;
            {4'd0, 3'd6, 3'd6}: kernel_rom_out = 16'sd13399;
            {4'd0, 3'd6, 3'd7}: kernel_rom_out = -16'sd8523;
            {4'd0, 3'd7, 3'd0}: kernel_rom_out = -16'sd10528;
            {4'd0, 3'd7, 3'd1}: kernel_rom_out = -16'sd12809;
            {4'd0, 3'd7, 3'd2}: kernel_rom_out = -16'sd11788;
            {4'd0, 3'd7, 3'd3}: kernel_rom_out = 16'sd12520;
            {4'd0, 3'd7, 3'd4}: kernel_rom_out = 16'sd14036;
            {4'd0, 3'd7, 3'd5}: kernel_rom_out = 16'sd14281;
            {4'd0, 3'd7, 3'd6}: kernel_rom_out = -16'sd9488;
            {4'd0, 3'd7, 3'd7}: kernel_rom_out = 16'sd3470;

            // MODE 1: RFT-FIBONACCI (unitarity: 1.09e-13)
            {4'd1, 3'd0, 3'd0}: kernel_rom_out = 16'sd3859;
            {4'd1, 3'd0, 3'd1}: kernel_rom_out = -16'sd9620;
            {4'd1, 3'd0, 3'd2}: kernel_rom_out = 16'sd15561;
            {4'd1, 3'd0, 3'd3}: kernel_rom_out = -16'sd13362;
            {4'd1, 3'd0, 3'd4}: kernel_rom_out = 16'sd11981;
            {4'd1, 3'd0, 3'd5}: kernel_rom_out = -16'sd11555;
            {4'd1, 3'd0, 3'd6}: kernel_rom_out = 16'sd11672;
            {4'd1, 3'd0, 3'd7}: kernel_rom_out = 16'sd11499;
            {4'd1, 3'd1, 3'd0}: kernel_rom_out = 16'sd8362;
            {4'd1, 3'd1, 3'd1}: kernel_rom_out = -16'sd13352;
            {4'd1, 3'd1, 3'd2}: kernel_rom_out = 16'sd14810;
            {4'd1, 3'd1, 3'd3}: kernel_rom_out = 16'sd9564;
            {4'd1, 3'd1, 3'd4}: kernel_rom_out = -16'sd10614;
            {4'd1, 3'd1, 3'd5}: kernel_rom_out = -16'sd11499;
            {4'd1, 3'd1, 3'd6}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd1, 3'd7}: kernel_rom_out = -16'sd11613;
            {4'd1, 3'd2, 3'd0}: kernel_rom_out = 16'sd12646;
            {4'd1, 3'd2, 3'd1}: kernel_rom_out = -16'sd13286;
            {4'd1, 3'd2, 3'd2}: kernel_rom_out = -16'sd5722;
            {4'd1, 3'd2, 3'd3}: kernel_rom_out = 16'sd9516;
            {4'd1, 3'd2, 3'd4}: kernel_rom_out = 16'sd14559;
            {4'd1, 3'd2, 3'd5}: kernel_rom_out = 16'sd11614;
            {4'd1, 3'd2, 3'd6}: kernel_rom_out = -16'sd11497;
            {4'd1, 3'd2, 3'd7}: kernel_rom_out = 16'sd11613;
            {4'd1, 3'd3, 3'd0}: kernel_rom_out = 16'sd17090;
            {4'd1, 3'd3, 3'd1}: kernel_rom_out = -16'sd9460;
            {4'd1, 3'd3, 3'd2}: kernel_rom_out = -16'sd6526;
            {4'd1, 3'd3, 3'd3}: kernel_rom_out = -16'sd13276;
            {4'd1, 3'd3, 3'd4}: kernel_rom_out = -16'sd8285;
            {4'd1, 3'd3, 3'd5}: kernel_rom_out = 16'sd11671;
            {4'd1, 3'd3, 3'd6}: kernel_rom_out = 16'sd11555;
            {4'd1, 3'd3, 3'd7}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd4, 3'd0}: kernel_rom_out = 16'sd17090;
            {4'd1, 3'd4, 3'd1}: kernel_rom_out = 16'sd9460;
            {4'd1, 3'd4, 3'd2}: kernel_rom_out = -16'sd6526;
            {4'd1, 3'd4, 3'd3}: kernel_rom_out = 16'sd13276;
            {4'd1, 3'd4, 3'd4}: kernel_rom_out = -16'sd8285;
            {4'd1, 3'd4, 3'd5}: kernel_rom_out = -16'sd11671;
            {4'd1, 3'd4, 3'd6}: kernel_rom_out = 16'sd11555;
            {4'd1, 3'd4, 3'd7}: kernel_rom_out = 16'sd11614;
            {4'd1, 3'd5, 3'd0}: kernel_rom_out = 16'sd12646;
            {4'd1, 3'd5, 3'd1}: kernel_rom_out = 16'sd13286;
            {4'd1, 3'd5, 3'd2}: kernel_rom_out = -16'sd5722;
            {4'd1, 3'd5, 3'd3}: kernel_rom_out = -16'sd9516;
            {4'd1, 3'd5, 3'd4}: kernel_rom_out = 16'sd14559;
            {4'd1, 3'd5, 3'd5}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd5, 3'd6}: kernel_rom_out = -16'sd11497;
            {4'd1, 3'd5, 3'd7}: kernel_rom_out = -16'sd11613;
            {4'd1, 3'd6, 3'd0}: kernel_rom_out = 16'sd8362;
            {4'd1, 3'd6, 3'd1}: kernel_rom_out = 16'sd13352;
            {4'd1, 3'd6, 3'd2}: kernel_rom_out = 16'sd14810;
            {4'd1, 3'd6, 3'd3}: kernel_rom_out = -16'sd9564;
            {4'd1, 3'd6, 3'd4}: kernel_rom_out = -16'sd10614;
            {4'd1, 3'd6, 3'd5}: kernel_rom_out = 16'sd11499;
            {4'd1, 3'd6, 3'd6}: kernel_rom_out = -16'sd11614;
            {4'd1, 3'd6, 3'd7}: kernel_rom_out = 16'sd11613;
            {4'd1, 3'd7, 3'd0}: kernel_rom_out = 16'sd3859;
            {4'd1, 3'd7, 3'd1}: kernel_rom_out = 16'sd9620;
            {4'd1, 3'd7, 3'd2}: kernel_rom_out = 16'sd15561;
            {4'd1, 3'd7, 3'd3}: kernel_rom_out = 16'sd13362;
            {4'd1, 3'd7, 3'd4}: kernel_rom_out = 16'sd11981;
            {4'd1, 3'd7, 3'd5}: kernel_rom_out = 16'sd11555;
            {4'd1, 3'd7, 3'd6}: kernel_rom_out = 16'sd11672;
            {4'd1, 3'd7, 3'd7}: kernel_rom_out = -16'sd11499;

            // MODE 2: RFT-HARMONIC (unitarity: 1.96e-15)
            {4'd2, 3'd0, 3'd0}: kernel_rom_out = 16'sd11505;
            {4'd2, 3'd0, 3'd1}: kernel_rom_out = -16'sd11573;
            {4'd2, 3'd0, 3'd2}: kernel_rom_out = 16'sd14539;
            {4'd2, 3'd0, 3'd3}: kernel_rom_out = 16'sd16484;
            {4'd2, 3'd0, 3'd4}: kernel_rom_out = 16'sd8842;
            {4'd2, 3'd0, 3'd5}: kernel_rom_out = -16'sd13592;
            {4'd2, 3'd0, 3'd6}: kernel_rom_out = 16'sd2596;
            {4'd2, 3'd0, 3'd7}: kernel_rom_out = 16'sd7386;
            {4'd2, 3'd1, 3'd0}: kernel_rom_out = -16'sd11549;
            {4'd2, 3'd1, 3'd1}: kernel_rom_out = -16'sd11481;
            {4'd2, 3'd1, 3'd2}: kernel_rom_out = -16'sd15661;
            {4'd2, 3'd1, 3'd3}: kernel_rom_out = 16'sd13444;
            {4'd2, 3'd1, 3'd4}: kernel_rom_out = -16'sd14106;
            {4'd2, 3'd1, 3'd5}: kernel_rom_out = -16'sd8723;
            {4'd2, 3'd1, 3'd6}: kernel_rom_out = -16'sd9147;
            {4'd2, 3'd1, 3'd7}: kernel_rom_out = 16'sd4871;
            {4'd2, 3'd2, 3'd0}: kernel_rom_out = 16'sd11635;
            {4'd2, 3'd2, 3'd1}: kernel_rom_out = -16'sd11657;
            {4'd2, 3'd2, 3'd2}: kernel_rom_out = 16'sd6800;
            {4'd2, 3'd2, 3'd3}: kernel_rom_out = 16'sd4852;
            {4'd2, 3'd2, 3'd4}: kernel_rom_out = -16'sd10542;
            {4'd2, 3'd2, 3'd5}: kernel_rom_out = 16'sd15032;
            {4'd2, 3'd2, 3'd6}: kernel_rom_out = -16'sd11345;
            {4'd2, 3'd2, 3'd7}: kernel_rom_out = -16'sd16334;
            {4'd2, 3'd3, 3'd0}: kernel_rom_out = -16'sd11649;
            {4'd2, 3'd3, 3'd1}: kernel_rom_out = -16'sd11626;
            {4'd2, 3'd3, 3'd2}: kernel_rom_out = -16'sd5826;
            {4'd2, 3'd3, 3'd3}: kernel_rom_out = 16'sd7797;
            {4'd2, 3'd3, 3'd4}: kernel_rom_out = 16'sd12188;
            {4'd2, 3'd3, 3'd5}: kernel_rom_out = 16'sd7072;
            {4'd2, 3'd3, 3'd6}: kernel_rom_out = 16'sd17824;
            {4'd2, 3'd3, 3'd7}: kernel_rom_out = -16'sd13848;
            {4'd2, 3'd4, 3'd0}: kernel_rom_out = 16'sd11649;
            {4'd2, 3'd4, 3'd1}: kernel_rom_out = -16'sd11626;
            {4'd2, 3'd4, 3'd2}: kernel_rom_out = -16'sd5826;
            {4'd2, 3'd4, 3'd3}: kernel_rom_out = -16'sd7797;
            {4'd2, 3'd4, 3'd4}: kernel_rom_out = -16'sd12188;
            {4'd2, 3'd4, 3'd5}: kernel_rom_out = 16'sd7072;
            {4'd2, 3'd4, 3'd6}: kernel_rom_out = 16'sd17824;
            {4'd2, 3'd4, 3'd7}: kernel_rom_out = 16'sd13848;
            {4'd2, 3'd5, 3'd0}: kernel_rom_out = -16'sd11635;
            {4'd2, 3'd5, 3'd1}: kernel_rom_out = -16'sd11657;
            {4'd2, 3'd5, 3'd2}: kernel_rom_out = 16'sd6800;
            {4'd2, 3'd5, 3'd3}: kernel_rom_out = -16'sd4852;
            {4'd2, 3'd5, 3'd4}: kernel_rom_out = 16'sd10542;
            {4'd2, 3'd5, 3'd5}: kernel_rom_out = 16'sd15032;
            {4'd2, 3'd5, 3'd6}: kernel_rom_out = -16'sd11345;
            {4'd2, 3'd5, 3'd7}: kernel_rom_out = 16'sd16334;
            {4'd2, 3'd6, 3'd0}: kernel_rom_out = 16'sd11549;
            {4'd2, 3'd6, 3'd1}: kernel_rom_out = -16'sd11481;
            {4'd2, 3'd6, 3'd2}: kernel_rom_out = -16'sd15661;
            {4'd2, 3'd6, 3'd3}: kernel_rom_out = -16'sd13444;
            {4'd2, 3'd6, 3'd4}: kernel_rom_out = 16'sd14106;
            {4'd2, 3'd6, 3'd5}: kernel_rom_out = -16'sd8723;
            {4'd2, 3'd6, 3'd6}: kernel_rom_out = -16'sd9147;
            {4'd2, 3'd6, 3'd7}: kernel_rom_out = -16'sd4871;
            {4'd2, 3'd7, 3'd0}: kernel_rom_out = -16'sd11505;
            {4'd2, 3'd7, 3'd1}: kernel_rom_out = -16'sd11573;
            {4'd2, 3'd7, 3'd2}: kernel_rom_out = 16'sd14539;
            {4'd2, 3'd7, 3'd3}: kernel_rom_out = -16'sd16484;
            {4'd2, 3'd7, 3'd4}: kernel_rom_out = -16'sd8842;
            {4'd2, 3'd7, 3'd5}: kernel_rom_out = -16'sd13592;
            {4'd2, 3'd7, 3'd6}: kernel_rom_out = 16'sd2596;
            {4'd2, 3'd7, 3'd7}: kernel_rom_out = -16'sd7386;

            // MODE 3: RFT-GEOMETRIC (unitarity: 3.58e-15)
            {4'd3, 3'd0, 3'd0}: kernel_rom_out = -16'sd13692;
            {4'd3, 3'd0, 3'd1}: kernel_rom_out = 16'sd663;
            {4'd3, 3'd0, 3'd2}: kernel_rom_out = 16'sd20505;
            {4'd3, 3'd0, 3'd3}: kernel_rom_out = -16'sd9236;
            {4'd3, 3'd0, 3'd4}: kernel_rom_out = -16'sd9709;
            {4'd3, 3'd0, 3'd5}: kernel_rom_out = -16'sd3379;
            {4'd3, 3'd0, 3'd6}: kernel_rom_out = 16'sd15895;
            {4'd3, 3'd0, 3'd7}: kernel_rom_out = -16'sd4653;
            {4'd3, 3'd1, 3'd0}: kernel_rom_out = -16'sd10201;
            {4'd3, 3'd1, 3'd1}: kernel_rom_out = 16'sd13503;
            {4'd3, 3'd1, 3'd2}: kernel_rom_out = 16'sd8329;
            {4'd3, 3'd1, 3'd3}: kernel_rom_out = 16'sd4498;
            {4'd3, 3'd1, 3'd4}: kernel_rom_out = 16'sd13956;
            {4'd3, 3'd1, 3'd5}: kernel_rom_out = 16'sd20225;
            {4'd3, 3'd1, 3'd6}: kernel_rom_out = -16'sd1874;
            {4'd3, 3'd1, 3'd7}: kernel_rom_out = 16'sd9506;
            {4'd3, 3'd2, 3'd0}: kernel_rom_out = 16'sd4467;
            {4'd3, 3'd2, 3'd1}: kernel_rom_out = 16'sd17252;
            {4'd3, 3'd2, 3'd2}: kernel_rom_out = -16'sd5562;
            {4'd3, 3'd2, 3'd3}: kernel_rom_out = 16'sd17817;
            {4'd3, 3'd2, 3'd4}: kernel_rom_out = -16'sd3910;
            {4'd3, 3'd2, 3'd5}: kernel_rom_out = -16'sd401;
            {4'd3, 3'd2, 3'd6}: kernel_rom_out = 16'sd14116;
            {4'd3, 3'd2, 3'd7}: kernel_rom_out = -16'sd13892;
            {4'd3, 3'd3, 3'd0}: kernel_rom_out = 16'sd15012;
            {4'd3, 3'd3, 3'd1}: kernel_rom_out = 16'sd7512;
            {4'd3, 3'd3, 3'd2}: kernel_rom_out = -16'sd4007;
            {4'd3, 3'd3, 3'd3}: kernel_rom_out = -16'sd10670;
            {4'd3, 3'd3, 3'd4}: kernel_rom_out = -16'sd15248;
            {4'd3, 3'd3, 3'd5}: kernel_rom_out = 16'sd10781;
            {4'd3, 3'd3, 3'd6}: kernel_rom_out = 16'sd9023;
            {4'd3, 3'd3, 3'd7}: kernel_rom_out = 16'sd15226;
            {4'd3, 3'd4, 3'd0}: kernel_rom_out = 16'sd15012;
            {4'd3, 3'd4, 3'd1}: kernel_rom_out = -16'sd7512;
            {4'd3, 3'd4, 3'd2}: kernel_rom_out = 16'sd4007;
            {4'd3, 3'd4, 3'd3}: kernel_rom_out = -16'sd10670;
            {4'd3, 3'd4, 3'd4}: kernel_rom_out = 16'sd15248;
            {4'd3, 3'd4, 3'd5}: kernel_rom_out = 16'sd10781;
            {4'd3, 3'd4, 3'd6}: kernel_rom_out = 16'sd9023;
            {4'd3, 3'd4, 3'd7}: kernel_rom_out = -16'sd15226;
            {4'd3, 3'd5, 3'd0}: kernel_rom_out = 16'sd4467;
            {4'd3, 3'd5, 3'd1}: kernel_rom_out = -16'sd17252;
            {4'd3, 3'd5, 3'd2}: kernel_rom_out = 16'sd5562;
            {4'd3, 3'd5, 3'd3}: kernel_rom_out = 16'sd17817;
            {4'd3, 3'd5, 3'd4}: kernel_rom_out = 16'sd3910;
            {4'd3, 3'd5, 3'd5}: kernel_rom_out = -16'sd401;
            {4'd3, 3'd5, 3'd6}: kernel_rom_out = 16'sd14116;
            {4'd3, 3'd5, 3'd7}: kernel_rom_out = 16'sd13892;
            {4'd3, 3'd6, 3'd0}: kernel_rom_out = -16'sd10201;
            {4'd3, 3'd6, 3'd1}: kernel_rom_out = -16'sd13503;
            {4'd3, 3'd6, 3'd2}: kernel_rom_out = -16'sd8329;
            {4'd3, 3'd6, 3'd3}: kernel_rom_out = 16'sd4498;
            {4'd3, 3'd6, 3'd4}: kernel_rom_out = -16'sd13956;
            {4'd3, 3'd6, 3'd5}: kernel_rom_out = 16'sd20225;
            {4'd3, 3'd6, 3'd6}: kernel_rom_out = -16'sd1874;
            {4'd3, 3'd6, 3'd7}: kernel_rom_out = -16'sd9506;
            {4'd3, 3'd7, 3'd0}: kernel_rom_out = -16'sd13692;
            {4'd3, 3'd7, 3'd1}: kernel_rom_out = -16'sd663;
            {4'd3, 3'd7, 3'd2}: kernel_rom_out = -16'sd20505;
            {4'd3, 3'd7, 3'd3}: kernel_rom_out = -16'sd9236;
            {4'd3, 3'd7, 3'd4}: kernel_rom_out = 16'sd9709;
            {4'd3, 3'd7, 3'd5}: kernel_rom_out = -16'sd3379;
            {4'd3, 3'd7, 3'd6}: kernel_rom_out = 16'sd15895;
            {4'd3, 3'd7, 3'd7}: kernel_rom_out = 16'sd4653;

            // MODE 4: RFT-BEATING (unitarity: 3.09e-15)
            {4'd4, 3'd0, 3'd0}: kernel_rom_out = -16'sd11094;
            {4'd4, 3'd0, 3'd1}: kernel_rom_out = 16'sd15417;
            {4'd4, 3'd0, 3'd2}: kernel_rom_out = 16'sd5892;
            {4'd4, 3'd0, 3'd3}: kernel_rom_out = -16'sd12981;
            {4'd4, 3'd0, 3'd4}: kernel_rom_out = 16'sd18457;
            {4'd4, 3'd0, 3'd5}: kernel_rom_out = -16'sd6279;
            {4'd4, 3'd0, 3'd6}: kernel_rom_out = 16'sd6194;
            {4'd4, 3'd0, 3'd7}: kernel_rom_out = -16'sd9551;
            {4'd4, 3'd1, 3'd0}: kernel_rom_out = -16'sd12220;
            {4'd4, 3'd1, 3'd1}: kernel_rom_out = -16'sd6858;
            {4'd4, 3'd1, 3'd2}: kernel_rom_out = -16'sd14172;
            {4'd4, 3'd1, 3'd3}: kernel_rom_out = -16'sd16386;
            {4'd4, 3'd1, 3'd4}: kernel_rom_out = -16'sd6798;
            {4'd4, 3'd1, 3'd5}: kernel_rom_out = 16'sd14804;
            {4'd4, 3'd1, 3'd6}: kernel_rom_out = 16'sd11852;
            {4'd4, 3'd1, 3'd7}: kernel_rom_out = 16'sd1466;
            {4'd4, 3'd2, 3'd0}: kernel_rom_out = -16'sd10860;
            {4'd4, 3'd2, 3'd1}: kernel_rom_out = -16'sd5461;
            {4'd4, 3'd2, 3'd2}: kernel_rom_out = 16'sd16367;
            {4'd4, 3'd2, 3'd3}: kernel_rom_out = -16'sd9717;
            {4'd4, 3'd2, 3'd4}: kernel_rom_out = -16'sd12212;
            {4'd4, 3'd2, 3'd5}: kernel_rom_out = -16'sd14677;
            {4'd4, 3'd2, 3'd6}: kernel_rom_out = 16'sd1369;
            {4'd4, 3'd2, 3'd7}: kernel_rom_out = 16'sd14042;
            {4'd4, 3'd3, 3'd0}: kernel_rom_out = -16'sd12104;
            {4'd4, 3'd3, 3'd1}: kernel_rom_out = 16'sd14909;
            {4'd4, 3'd3, 3'd2}: kernel_rom_out = -16'sd5778;
            {4'd4, 3'd3, 3'd3}: kernel_rom_out = 16'sd2326;
            {4'd4, 3'd3, 3'd4}: kernel_rom_out = 16'sd903;
            {4'd4, 3'd3, 3'd5}: kernel_rom_out = 16'sd7927;
            {4'd4, 3'd3, 3'd6}: kernel_rom_out = -16'sd18871;
            {4'd4, 3'd3, 3'd7}: kernel_rom_out = 16'sd15694;
            {4'd4, 3'd4, 3'd0}: kernel_rom_out = -16'sd12104;
            {4'd4, 3'd4, 3'd1}: kernel_rom_out = -16'sd14909;
            {4'd4, 3'd4, 3'd2}: kernel_rom_out = -16'sd5778;
            {4'd4, 3'd4, 3'd3}: kernel_rom_out = -16'sd2326;
            {4'd4, 3'd4, 3'd4}: kernel_rom_out = 16'sd903;
            {4'd4, 3'd4, 3'd5}: kernel_rom_out = -16'sd7927;
            {4'd4, 3'd4, 3'd6}: kernel_rom_out = -16'sd18871;
            {4'd4, 3'd4, 3'd7}: kernel_rom_out = -16'sd15694;
            {4'd4, 3'd5, 3'd0}: kernel_rom_out = -16'sd10860;
            {4'd4, 3'd5, 3'd1}: kernel_rom_out = 16'sd5461;
            {4'd4, 3'd5, 3'd2}: kernel_rom_out = 16'sd16367;
            {4'd4, 3'd5, 3'd3}: kernel_rom_out = 16'sd9717;
            {4'd4, 3'd5, 3'd4}: kernel_rom_out = -16'sd12212;
            {4'd4, 3'd5, 3'd5}: kernel_rom_out = 16'sd14677;
            {4'd4, 3'd5, 3'd6}: kernel_rom_out = 16'sd1369;
            {4'd4, 3'd5, 3'd7}: kernel_rom_out = -16'sd14042;
            {4'd4, 3'd6, 3'd0}: kernel_rom_out = -16'sd12220;
            {4'd4, 3'd6, 3'd1}: kernel_rom_out = 16'sd6858;
            {4'd4, 3'd6, 3'd2}: kernel_rom_out = -16'sd14172;
            {4'd4, 3'd6, 3'd3}: kernel_rom_out = 16'sd16386;
            {4'd4, 3'd6, 3'd4}: kernel_rom_out = -16'sd6798;
            {4'd4, 3'd6, 3'd5}: kernel_rom_out = -16'sd14804;
            {4'd4, 3'd6, 3'd6}: kernel_rom_out = 16'sd11852;
            {4'd4, 3'd6, 3'd7}: kernel_rom_out = -16'sd1466;
            {4'd4, 3'd7, 3'd0}: kernel_rom_out = -16'sd11094;
            {4'd4, 3'd7, 3'd1}: kernel_rom_out = -16'sd15417;
            {4'd4, 3'd7, 3'd2}: kernel_rom_out = 16'sd5892;
            {4'd4, 3'd7, 3'd3}: kernel_rom_out = 16'sd12981;
            {4'd4, 3'd7, 3'd4}: kernel_rom_out = 16'sd18457;
            {4'd4, 3'd7, 3'd5}: kernel_rom_out = 16'sd6279;
            {4'd4, 3'd7, 3'd6}: kernel_rom_out = 16'sd6194;
            {4'd4, 3'd7, 3'd7}: kernel_rom_out = 16'sd9551;

            // MODE 5: RFT-PHYLLOTAXIS (unitarity: 4.38e-15)
            {4'd5, 3'd0, 3'd0}: kernel_rom_out = 16'sd9597;
            {4'd5, 3'd0, 3'd1}: kernel_rom_out = 16'sd15505;
            {4'd5, 3'd0, 3'd2}: kernel_rom_out = -16'sd9608;
            {4'd5, 3'd0, 3'd3}: kernel_rom_out = 16'sd5574;
            {4'd5, 3'd0, 3'd4}: kernel_rom_out = 16'sd13824;
            {4'd5, 3'd0, 3'd5}: kernel_rom_out = -16'sd3604;
            {4'd5, 3'd0, 3'd6}: kernel_rom_out = 16'sd16222;
            {4'd5, 3'd0, 3'd7}: kernel_rom_out = -16'sd12268;
            {4'd5, 3'd1, 3'd0}: kernel_rom_out = -16'sd16171;
            {4'd5, 3'd1, 3'd1}: kernel_rom_out = -16'sd1835;
            {4'd5, 3'd1, 3'd2}: kernel_rom_out = 16'sd248;
            {4'd5, 3'd1, 3'd3}: kernel_rom_out = 16'sd12282;
            {4'd5, 3'd1, 3'd4}: kernel_rom_out = 16'sd7890;
            {4'd5, 3'd1, 3'd5}: kernel_rom_out = 16'sd21706;
            {4'd5, 3'd1, 3'd6}: kernel_rom_out = -16'sd2818;
            {4'd5, 3'd1, 3'd7}: kernel_rom_out = -16'sd10796;
            {4'd5, 3'd2, 3'd0}: kernel_rom_out = 16'sd12685;
            {4'd5, 3'd2, 3'd1}: kernel_rom_out = -16'sd11019;
            {4'd5, 3'd2, 3'd2}: kernel_rom_out = 16'sd9066;
            {4'd5, 3'd2, 3'd3}: kernel_rom_out = 16'sd4638;
            {4'd5, 3'd2, 3'd4}: kernel_rom_out = 16'sd16799;
            {4'd5, 3'd2, 3'd5}: kernel_rom_out = -16'sd7142;
            {4'd5, 3'd2, 3'd6}: kernel_rom_out = -16'sd16266;
            {4'd5, 3'd2, 3'd7}: kernel_rom_out = -16'sd9477;
            {4'd5, 3'd3, 3'd0}: kernel_rom_out = -16'sd4725;
            {4'd5, 3'd3, 3'd1}: kernel_rom_out = 16'sd13100;
            {4'd5, 3'd3, 3'd2}: kernel_rom_out = 16'sd19033;
            {4'd5, 3'd3, 3'd3}: kernel_rom_out = -16'sd18259;
            {4'd5, 3'd3, 3'd4}: kernel_rom_out = -16'sd1126;
            {4'd5, 3'd3, 3'd5}: kernel_rom_out = 16'sd1299;
            {4'd5, 3'd3, 3'd6}: kernel_rom_out = -16'sd1075;
            {4'd5, 3'd3, 3'd7}: kernel_rom_out = -16'sd13415;
            {4'd5, 3'd4, 3'd0}: kernel_rom_out = -16'sd4725;
            {4'd5, 3'd4, 3'd1}: kernel_rom_out = -16'sd13100;
            {4'd5, 3'd4, 3'd2}: kernel_rom_out = -16'sd19033;
            {4'd5, 3'd4, 3'd3}: kernel_rom_out = -16'sd18259;
            {4'd5, 3'd4, 3'd4}: kernel_rom_out = 16'sd1126;
            {4'd5, 3'd4, 3'd5}: kernel_rom_out = -16'sd1299;
            {4'd5, 3'd4, 3'd6}: kernel_rom_out = -16'sd1075;
            {4'd5, 3'd4, 3'd7}: kernel_rom_out = -16'sd13415;
            {4'd5, 3'd5, 3'd0}: kernel_rom_out = 16'sd12685;
            {4'd5, 3'd5, 3'd1}: kernel_rom_out = 16'sd11019;
            {4'd5, 3'd5, 3'd2}: kernel_rom_out = -16'sd9066;
            {4'd5, 3'd5, 3'd3}: kernel_rom_out = 16'sd4638;
            {4'd5, 3'd5, 3'd4}: kernel_rom_out = -16'sd16799;
            {4'd5, 3'd5, 3'd5}: kernel_rom_out = 16'sd7142;
            {4'd5, 3'd5, 3'd6}: kernel_rom_out = -16'sd16266;
            {4'd5, 3'd5, 3'd7}: kernel_rom_out = -16'sd9477;
            {4'd5, 3'd6, 3'd0}: kernel_rom_out = -16'sd16171;
            {4'd5, 3'd6, 3'd1}: kernel_rom_out = 16'sd1835;
            {4'd5, 3'd6, 3'd2}: kernel_rom_out = -16'sd248;
            {4'd5, 3'd6, 3'd3}: kernel_rom_out = 16'sd12282;
            {4'd5, 3'd6, 3'd4}: kernel_rom_out = -16'sd7890;
            {4'd5, 3'd6, 3'd5}: kernel_rom_out = -16'sd21706;
            {4'd5, 3'd6, 3'd6}: kernel_rom_out = -16'sd2818;
            {4'd5, 3'd6, 3'd7}: kernel_rom_out = -16'sd10796;
            {4'd5, 3'd7, 3'd0}: kernel_rom_out = 16'sd9597;
            {4'd5, 3'd7, 3'd1}: kernel_rom_out = -16'sd15505;
            {4'd5, 3'd7, 3'd2}: kernel_rom_out = 16'sd9608;
            {4'd5, 3'd7, 3'd3}: kernel_rom_out = 16'sd5574;
            {4'd5, 3'd7, 3'd4}: kernel_rom_out = -16'sd13824;
            {4'd5, 3'd7, 3'd5}: kernel_rom_out = 16'sd3604;
            {4'd5, 3'd7, 3'd6}: kernel_rom_out = 16'sd16222;
            {4'd5, 3'd7, 3'd7}: kernel_rom_out = -16'sd12268;

            // MODE 6: RFT-CASCADE (unitarity: 1.51e-15)
            {4'd6, 3'd0, 3'd0}: kernel_rom_out = -16'sd9727;
            {4'd6, 3'd0, 3'd1}: kernel_rom_out = 16'sd15910;
            {4'd6, 3'd0, 3'd2}: kernel_rom_out = 16'sd14164;
            {4'd6, 3'd0, 3'd3}: kernel_rom_out = -16'sd2527;
            {4'd6, 3'd0, 3'd4}: kernel_rom_out = 16'sd15410;
            {4'd6, 3'd0, 3'd5}: kernel_rom_out = -16'sd4311;
            {4'd6, 3'd0, 3'd6}: kernel_rom_out = 16'sd2029;
            {4'd6, 3'd0, 3'd7}: kernel_rom_out = 16'sd16085;
            {4'd6, 3'd1, 3'd0}: kernel_rom_out = -16'sd10888;
            {4'd6, 3'd1, 3'd1}: kernel_rom_out = 16'sd16012;
            {4'd6, 3'd1, 3'd2}: kernel_rom_out = -16'sd12647;
            {4'd6, 3'd1, 3'd3}: kernel_rom_out = -16'sd3171;
            {4'd6, 3'd1, 3'd4}: kernel_rom_out = 16'sd2664;
            {4'd6, 3'd1, 3'd5}: kernel_rom_out = 16'sd8553;
            {4'd6, 3'd1, 3'd6}: kernel_rom_out = 16'sd15851;
            {4'd6, 3'd1, 3'd7}: kernel_rom_out = -16'sd14044;
            {4'd6, 3'd2, 3'd0}: kernel_rom_out = -16'sd12549;
            {4'd6, 3'd2, 3'd1}: kernel_rom_out = -16'sd1629;
            {4'd6, 3'd2, 3'd2}: kernel_rom_out = -16'sd9517;
            {4'd6, 3'd2, 3'd3}: kernel_rom_out = -16'sd19434;
            {4'd6, 3'd2, 3'd4}: kernel_rom_out = 16'sd3029;
            {4'd6, 3'd2, 3'd5}: kernel_rom_out = -16'sd11648;
            {4'd6, 3'd2, 3'd6}: kernel_rom_out = -16'sd16722;
            {4'd6, 3'd2, 3'd7}: kernel_rom_out = -16'sd4564;
            {4'd6, 3'd3, 3'd0}: kernel_rom_out = -16'sd12892;
            {4'd6, 3'd3, 3'd1}: kernel_rom_out = -16'sd4965;
            {4'd6, 3'd3, 3'd2}: kernel_rom_out = 16'sd9257;
            {4'd6, 3'd3, 3'd3}: kernel_rom_out = -16'sd11946;
            {4'd6, 3'd3, 3'd4}: kernel_rom_out = -16'sd16825;
            {4'd6, 3'd3, 3'd5}: kernel_rom_out = 16'sd17590;
            {4'd6, 3'd3, 3'd6}: kernel_rom_out = 16'sd1358;
            {4'd6, 3'd3, 3'd7}: kernel_rom_out = 16'sd7749;
            {4'd6, 3'd4, 3'd0}: kernel_rom_out = -16'sd12892;
            {4'd6, 3'd4, 3'd1}: kernel_rom_out = 16'sd4965;
            {4'd6, 3'd4, 3'd2}: kernel_rom_out = 16'sd9257;
            {4'd6, 3'd4, 3'd3}: kernel_rom_out = 16'sd11946;
            {4'd6, 3'd4, 3'd4}: kernel_rom_out = -16'sd16825;
            {4'd6, 3'd4, 3'd5}: kernel_rom_out = -16'sd17590;
            {4'd6, 3'd4, 3'd6}: kernel_rom_out = 16'sd1358;
            {4'd6, 3'd4, 3'd7}: kernel_rom_out = -16'sd7749;
            {4'd6, 3'd5, 3'd0}: kernel_rom_out = -16'sd12549;
            {4'd6, 3'd5, 3'd1}: kernel_rom_out = 16'sd1629;
            {4'd6, 3'd5, 3'd2}: kernel_rom_out = -16'sd9517;
            {4'd6, 3'd5, 3'd3}: kernel_rom_out = 16'sd19434;
            {4'd6, 3'd5, 3'd4}: kernel_rom_out = 16'sd3029;
            {4'd6, 3'd5, 3'd5}: kernel_rom_out = 16'sd11648;
            {4'd6, 3'd5, 3'd6}: kernel_rom_out = -16'sd16722;
            {4'd6, 3'd5, 3'd7}: kernel_rom_out = 16'sd4564;
            {4'd6, 3'd6, 3'd0}: kernel_rom_out = -16'sd10888;
            {4'd6, 3'd6, 3'd1}: kernel_rom_out = -16'sd16012;
            {4'd6, 3'd6, 3'd2}: kernel_rom_out = -16'sd12647;
            {4'd6, 3'd6, 3'd3}: kernel_rom_out = 16'sd3171;
            {4'd6, 3'd6, 3'd4}: kernel_rom_out = 16'sd2664;
            {4'd6, 3'd6, 3'd5}: kernel_rom_out = -16'sd8553;
            {4'd6, 3'd6, 3'd6}: kernel_rom_out = 16'sd15851;
            {4'd6, 3'd6, 3'd7}: kernel_rom_out = 16'sd14044;
            {4'd6, 3'd7, 3'd0}: kernel_rom_out = -16'sd9727;
            {4'd6, 3'd7, 3'd1}: kernel_rom_out = -16'sd15910;
            {4'd6, 3'd7, 3'd2}: kernel_rom_out = 16'sd14164;
            {4'd6, 3'd7, 3'd3}: kernel_rom_out = 16'sd2527;
            {4'd6, 3'd7, 3'd4}: kernel_rom_out = 16'sd15410;
            {4'd6, 3'd7, 3'd5}: kernel_rom_out = 16'sd4311;
            {4'd6, 3'd7, 3'd6}: kernel_rom_out = 16'sd2029;
            {4'd6, 3'd7, 3'd7}: kernel_rom_out = -16'sd16085;

            // MODE 7: RFT-HYBRID_DCT (unitarity: 1.12e-15)
            {4'd7, 3'd0, 3'd0}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd1}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd2}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd3}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd4}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd5}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd6}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd0, 3'd7}: kernel_rom_out = -16'sd11585;
            {4'd7, 3'd1, 3'd0}: kernel_rom_out = -16'sd16069;
            {4'd7, 3'd1, 3'd1}: kernel_rom_out = -16'sd13622;
            {4'd7, 3'd1, 3'd2}: kernel_rom_out = -16'sd9102;
            {4'd7, 3'd1, 3'd3}: kernel_rom_out = -16'sd3196;
            {4'd7, 3'd1, 3'd4}: kernel_rom_out = 16'sd3196;
            {4'd7, 3'd1, 3'd5}: kernel_rom_out = 16'sd9102;
            {4'd7, 3'd1, 3'd6}: kernel_rom_out = 16'sd13622;
            {4'd7, 3'd1, 3'd7}: kernel_rom_out = 16'sd16069;
            {4'd7, 3'd2, 3'd0}: kernel_rom_out = 16'sd15136;
            {4'd7, 3'd2, 3'd1}: kernel_rom_out = 16'sd6269;
            {4'd7, 3'd2, 3'd2}: kernel_rom_out = -16'sd6269;
            {4'd7, 3'd2, 3'd3}: kernel_rom_out = -16'sd15136;
            {4'd7, 3'd2, 3'd4}: kernel_rom_out = -16'sd15136;
            {4'd7, 3'd2, 3'd5}: kernel_rom_out = -16'sd6269;
            {4'd7, 3'd2, 3'd6}: kernel_rom_out = 16'sd6269;
            {4'd7, 3'd2, 3'd7}: kernel_rom_out = 16'sd15136;
            {4'd7, 3'd3, 3'd0}: kernel_rom_out = 16'sd13622;
            {4'd7, 3'd3, 3'd1}: kernel_rom_out = -16'sd3196;
            {4'd7, 3'd3, 3'd2}: kernel_rom_out = -16'sd16069;
            {4'd7, 3'd3, 3'd3}: kernel_rom_out = -16'sd9102;
            {4'd7, 3'd3, 3'd4}: kernel_rom_out = 16'sd9102;
            {4'd7, 3'd3, 3'd5}: kernel_rom_out = 16'sd16069;
            {4'd7, 3'd3, 3'd6}: kernel_rom_out = 16'sd3196;
            {4'd7, 3'd3, 3'd7}: kernel_rom_out = -16'sd13622;
            {4'd7, 3'd4, 3'd0}: kernel_rom_out = -16'sd9051;
            {4'd7, 3'd4, 3'd1}: kernel_rom_out = 16'sd15560;
            {4'd7, 3'd4, 3'd2}: kernel_rom_out = -16'sd9371;
            {4'd7, 3'd4, 3'd3}: kernel_rom_out = 16'sd10393;
            {4'd7, 3'd4, 3'd4}: kernel_rom_out = -16'sd15759;
            {4'd7, 3'd4, 3'd5}: kernel_rom_out = 16'sd4982;
            {4'd7, 3'd4, 3'd6}: kernel_rom_out = 16'sd13356;
            {4'd7, 3'd4, 3'd7}: kernel_rom_out = -16'sd10111;
            {4'd7, 3'd5, 3'd0}: kernel_rom_out = 16'sd2248;
            {4'd7, 3'd5, 3'd1}: kernel_rom_out = -16'sd7751;
            {4'd7, 3'd5, 3'd2}: kernel_rom_out = 16'sd10583;
            {4'd7, 3'd5, 3'd3}: kernel_rom_out = -16'sd6173;
            {4'd7, 3'd5, 3'd4}: kernel_rom_out = 16'sd3647;
            {4'd7, 3'd5, 3'd5}: kernel_rom_out = -16'sd13262;
            {4'd7, 3'd5, 3'd6}: kernel_rom_out = 16'sd22846;
            {4'd7, 3'd5, 3'd7}: kernel_rom_out = -16'sd12137;
            {4'd7, 3'd6, 3'd0}: kernel_rom_out = -16'sd7156;
            {4'd7, 3'd6, 3'd1}: kernel_rom_out = 16'sd3009;
            {4'd7, 3'd6, 3'd2}: kernel_rom_out = 16'sd18306;
            {4'd7, 3'd6, 3'd3}: kernel_rom_out = -16'sd16873;
            {4'd7, 3'd6, 3'd4}: kernel_rom_out = -16'sd8604;
            {4'd7, 3'd6, 3'd5}: kernel_rom_out = 16'sd17310;
            {4'd7, 3'd6, 3'd6}: kernel_rom_out = -16'sd2008;
            {4'd7, 3'd6, 3'd7}: kernel_rom_out = -16'sd3983;
            {4'd7, 3'd7, 3'd0}: kernel_rom_out = -16'sd11331;
            {4'd7, 3'd7, 3'd1}: kernel_rom_out = 16'sd19827;
            {4'd7, 3'd7, 3'd2}: kernel_rom_out = -16'sd4917;
            {4'd7, 3'd7, 3'd3}: kernel_rom_out = -16'sd13655;
            {4'd7, 3'd7, 3'd4}: kernel_rom_out = 16'sd16781;
            {4'd7, 3'd7, 3'd5}: kernel_rom_out = -16'sd7665;
            {4'd7, 3'd7, 3'd6}: kernel_rom_out = -16'sd122;
            {4'd7, 3'd7, 3'd7}: kernel_rom_out = 16'sd1083;

            // MODE 8: RFT-MANIFOLD (unitarity: 2.26e-15)
            {4'd8, 3'd0, 3'd0}: kernel_rom_out = -16'sd9374;
            {4'd8, 3'd0, 3'd1}: kernel_rom_out = -16'sd14997;
            {4'd8, 3'd0, 3'd2}: kernel_rom_out = -16'sd10409;
            {4'd8, 3'd0, 3'd3}: kernel_rom_out = -16'sd14601;
            {4'd8, 3'd0, 3'd4}: kernel_rom_out = -16'sd2148;
            {4'd8, 3'd0, 3'd5}: kernel_rom_out = -16'sd6335;
            {4'd8, 3'd0, 3'd6}: kernel_rom_out = -16'sd7654;
            {4'd8, 3'd0, 3'd7}: kernel_rom_out = 16'sd18330;
            {4'd8, 3'd1, 3'd0}: kernel_rom_out = -16'sd15451;
            {4'd8, 3'd1, 3'd1}: kernel_rom_out = -16'sd2699;
            {4'd8, 3'd1, 3'd2}: kernel_rom_out = 16'sd14530;
            {4'd8, 3'd1, 3'd3}: kernel_rom_out = -16'sd4158;
            {4'd8, 3'd1, 3'd4}: kernel_rom_out = 16'sd9216;
            {4'd8, 3'd1, 3'd5}: kernel_rom_out = -16'sd9076;
            {4'd8, 3'd1, 3'd6}: kernel_rom_out = 16'sd20734;
            {4'd8, 3'd1, 3'd7}: kernel_rom_out = 16'sd1429;
            {4'd8, 3'd2, 3'd0}: kernel_rom_out = -16'sd13688;
            {4'd8, 3'd2, 3'd1}: kernel_rom_out = 16'sd9764;
            {4'd8, 3'd2, 3'd2}: kernel_rom_out = -16'sd12176;
            {4'd8, 3'd2, 3'd3}: kernel_rom_out = 16'sd2159;
            {4'd8, 3'd2, 3'd4}: kernel_rom_out = -16'sd1565;
            {4'd8, 3'd2, 3'd5}: kernel_rom_out = -16'sd19719;
            {4'd8, 3'd2, 3'd6}: kernel_rom_out = -16'sd6927;
            {4'd8, 3'd2, 3'd7}: kernel_rom_out = -16'sd14099;
            {4'd8, 3'd3, 3'd0}: kernel_rom_out = -16'sd4780;
            {4'd8, 3'd3, 3'd1}: kernel_rom_out = 16'sd14468;
            {4'd8, 3'd3, 3'd2}: kernel_rom_out = 16'sd8313;
            {4'd8, 3'd3, 3'd3}: kernel_rom_out = -16'sd17369;
            {4'd8, 3'd3, 3'd4}: kernel_rom_out = -16'sd21091;
            {4'd8, 3'd3, 3'd5}: kernel_rom_out = 16'sd5047;
            {4'd8, 3'd3, 3'd6}: kernel_rom_out = 16'sd609;
            {4'd8, 3'd3, 3'd7}: kernel_rom_out = -16'sd196;
            {4'd8, 3'd4, 3'd0}: kernel_rom_out = 16'sd4780;
            {4'd8, 3'd4, 3'd1}: kernel_rom_out = 16'sd14468;
            {4'd8, 3'd4, 3'd2}: kernel_rom_out = -16'sd8313;
            {4'd8, 3'd4, 3'd3}: kernel_rom_out = -16'sd17369;
            {4'd8, 3'd4, 3'd4}: kernel_rom_out = 16'sd21091;
            {4'd8, 3'd4, 3'd5}: kernel_rom_out = 16'sd5047;
            {4'd8, 3'd4, 3'd6}: kernel_rom_out = 16'sd609;
            {4'd8, 3'd4, 3'd7}: kernel_rom_out = 16'sd196;
            {4'd8, 3'd5, 3'd0}: kernel_rom_out = 16'sd13688;
            {4'd8, 3'd5, 3'd1}: kernel_rom_out = 16'sd9764;
            {4'd8, 3'd5, 3'd2}: kernel_rom_out = 16'sd12176;
            {4'd8, 3'd5, 3'd3}: kernel_rom_out = 16'sd2159;
            {4'd8, 3'd5, 3'd4}: kernel_rom_out = 16'sd1565;
            {4'd8, 3'd5, 3'd5}: kernel_rom_out = -16'sd19719;
            {4'd8, 3'd5, 3'd6}: kernel_rom_out = -16'sd6927;
            {4'd8, 3'd5, 3'd7}: kernel_rom_out = 16'sd14099;
            {4'd8, 3'd6, 3'd0}: kernel_rom_out = 16'sd15451;
            {4'd8, 3'd6, 3'd1}: kernel_rom_out = -16'sd2699;
            {4'd8, 3'd6, 3'd2}: kernel_rom_out = -16'sd14530;
            {4'd8, 3'd6, 3'd3}: kernel_rom_out = -16'sd4158;
            {4'd8, 3'd6, 3'd4}: kernel_rom_out = -16'sd9216;
            {4'd8, 3'd6, 3'd5}: kernel_rom_out = -16'sd9076;
            {4'd8, 3'd6, 3'd6}: kernel_rom_out = 16'sd20734;
            {4'd8, 3'd6, 3'd7}: kernel_rom_out = -16'sd1429;
            {4'd8, 3'd7, 3'd0}: kernel_rom_out = 16'sd9374;
            {4'd8, 3'd7, 3'd1}: kernel_rom_out = -16'sd14997;
            {4'd8, 3'd7, 3'd2}: kernel_rom_out = 16'sd10409;
            {4'd8, 3'd7, 3'd3}: kernel_rom_out = -16'sd14601;
            {4'd8, 3'd7, 3'd4}: kernel_rom_out = 16'sd2148;
            {4'd8, 3'd7, 3'd5}: kernel_rom_out = -16'sd6335;
            {4'd8, 3'd7, 3'd6}: kernel_rom_out = -16'sd7654;
            {4'd8, 3'd7, 3'd7}: kernel_rom_out = -16'sd18330;

            // MODE 9: RFT-EULER (unitarity: 3.02e-15)
            {4'd9, 3'd0, 3'd0}: kernel_rom_out = -16'sd16232;
            {4'd9, 3'd0, 3'd1}: kernel_rom_out = 16'sd5203;
            {4'd9, 3'd0, 3'd2}: kernel_rom_out = -16'sd3776;
            {4'd9, 3'd0, 3'd3}: kernel_rom_out = -16'sd11809;
            {4'd9, 3'd0, 3'd4}: kernel_rom_out = 16'sd19982;
            {4'd9, 3'd0, 3'd5}: kernel_rom_out = -16'sd4049;
            {4'd9, 3'd0, 3'd6}: kernel_rom_out = 16'sd9809;
            {4'd9, 3'd0, 3'd7}: kernel_rom_out = -16'sd10839;
            {4'd9, 3'd1, 3'd0}: kernel_rom_out = -16'sd2338;
            {4'd9, 3'd1, 3'd1}: kernel_rom_out = 16'sd18201;
            {4'd9, 3'd1, 3'd2}: kernel_rom_out = -16'sd5501;
            {4'd9, 3'd1, 3'd3}: kernel_rom_out = -16'sd14165;
            {4'd9, 3'd1, 3'd4}: kernel_rom_out = -16'sd10024;
            {4'd9, 3'd1, 3'd5}: kernel_rom_out = 16'sd9963;
            {4'd9, 3'd1, 3'd6}: kernel_rom_out = 16'sd8648;
            {4'd9, 3'd1, 3'd7}: kernel_rom_out = 16'sd15213;
            {4'd9, 3'd2, 3'd0}: kernel_rom_out = 16'sd13633;
            {4'd9, 3'd2, 3'd1}: kernel_rom_out = 16'sd7122;
            {4'd9, 3'd2, 3'd2}: kernel_rom_out = -16'sd12391;
            {4'd9, 3'd2, 3'd3}: kernel_rom_out = -16'sd13010;
            {4'd9, 3'd2, 3'd4}: kernel_rom_out = 16'sd4481;
            {4'd9, 3'd2, 3'd5}: kernel_rom_out = -16'sd13424;
            {4'd9, 3'd2, 3'd6}: kernel_rom_out = -16'sd17677;
            {4'd9, 3'd2, 3'd7}: kernel_rom_out = -16'sd1227;
            {4'd9, 3'd3, 3'd0}: kernel_rom_out = 16'sd9056;
            {4'd9, 3'd3, 3'd1}: kernel_rom_out = -16'sd11303;
            {4'd9, 3'd3, 3'd2}: kernel_rom_out = -16'sd18406;
            {4'd9, 3'd3, 3'd3}: kernel_rom_out = -16'sd5239;
            {4'd9, 3'd3, 3'd4}: kernel_rom_out = -16'sd4120;
            {4'd9, 3'd3, 3'd5}: kernel_rom_out = 16'sd15523;
            {4'd9, 3'd3, 3'd6}: kernel_rom_out = 16'sd7303;
            {4'd9, 3'd3, 3'd7}: kernel_rom_out = -16'sd13653;
            {4'd9, 3'd4, 3'd0}: kernel_rom_out = -16'sd9056;
            {4'd9, 3'd4, 3'd1}: kernel_rom_out = -16'sd11303;
            {4'd9, 3'd4, 3'd2}: kernel_rom_out = -16'sd18406;
            {4'd9, 3'd4, 3'd3}: kernel_rom_out = 16'sd5239;
            {4'd9, 3'd4, 3'd4}: kernel_rom_out = -16'sd4120;
            {4'd9, 3'd4, 3'd5}: kernel_rom_out = -16'sd15523;
            {4'd9, 3'd4, 3'd6}: kernel_rom_out = 16'sd7303;
            {4'd9, 3'd4, 3'd7}: kernel_rom_out = 16'sd13653;
            {4'd9, 3'd5, 3'd0}: kernel_rom_out = -16'sd13633;
            {4'd9, 3'd5, 3'd1}: kernel_rom_out = 16'sd7122;
            {4'd9, 3'd5, 3'd2}: kernel_rom_out = -16'sd12391;
            {4'd9, 3'd5, 3'd3}: kernel_rom_out = 16'sd13010;
            {4'd9, 3'd5, 3'd4}: kernel_rom_out = 16'sd4481;
            {4'd9, 3'd5, 3'd5}: kernel_rom_out = 16'sd13424;
            {4'd9, 3'd5, 3'd6}: kernel_rom_out = -16'sd17677;
            {4'd9, 3'd5, 3'd7}: kernel_rom_out = 16'sd1227;
            {4'd9, 3'd6, 3'd0}: kernel_rom_out = 16'sd2338;
            {4'd9, 3'd6, 3'd1}: kernel_rom_out = 16'sd18201;
            {4'd9, 3'd6, 3'd2}: kernel_rom_out = -16'sd5501;
            {4'd9, 3'd6, 3'd3}: kernel_rom_out = 16'sd14165;
            {4'd9, 3'd6, 3'd4}: kernel_rom_out = -16'sd10024;
            {4'd9, 3'd6, 3'd5}: kernel_rom_out = -16'sd9963;
            {4'd9, 3'd6, 3'd6}: kernel_rom_out = 16'sd8648;
            {4'd9, 3'd6, 3'd7}: kernel_rom_out = -16'sd15213;
            {4'd9, 3'd7, 3'd0}: kernel_rom_out = 16'sd16232;
            {4'd9, 3'd7, 3'd1}: kernel_rom_out = 16'sd5203;
            {4'd9, 3'd7, 3'd2}: kernel_rom_out = -16'sd3776;
            {4'd9, 3'd7, 3'd3}: kernel_rom_out = 16'sd11809;
            {4'd9, 3'd7, 3'd4}: kernel_rom_out = 16'sd19982;
            {4'd9, 3'd7, 3'd5}: kernel_rom_out = 16'sd4049;
            {4'd9, 3'd7, 3'd6}: kernel_rom_out = 16'sd9809;
            {4'd9, 3'd7, 3'd7}: kernel_rom_out = 16'sd10839;

            // MODE 10: RFT-PHASE_COH (unitarity: 3.36e-15)
            {4'd10, 3'd0, 3'd0}: kernel_rom_out = -16'sd11229;
            {4'd10, 3'd0, 3'd1}: kernel_rom_out = -16'sd15554;
            {4'd10, 3'd0, 3'd2}: kernel_rom_out = 16'sd5617;
            {4'd10, 3'd0, 3'd3}: kernel_rom_out = -16'sd13614;
            {4'd10, 3'd0, 3'd4}: kernel_rom_out = -16'sd14765;
            {4'd10, 3'd0, 3'd5}: kernel_rom_out = 16'sd2171;
            {4'd10, 3'd0, 3'd6}: kernel_rom_out = 16'sd10240;
            {4'd10, 3'd0, 3'd7}: kernel_rom_out = 16'sd12696;
            {4'd10, 3'd1, 3'd0}: kernel_rom_out = -16'sd11768;
            {4'd10, 3'd1, 3'd1}: kernel_rom_out = 16'sd6617;
            {4'd10, 3'd1, 3'd2}: kernel_rom_out = -16'sd14607;
            {4'd10, 3'd1, 3'd3}: kernel_rom_out = -16'sd16824;
            {4'd10, 3'd1, 3'd4}: kernel_rom_out = 16'sd10658;
            {4'd10, 3'd1, 3'd5}: kernel_rom_out = 16'sd5380;
            {4'd10, 3'd1, 3'd6}: kernel_rom_out = -16'sd13456;
            {4'd10, 3'd1, 3'd7}: kernel_rom_out = 16'sd8449;
            {4'd10, 3'd2, 3'd0}: kernel_rom_out = -16'sd11428;
            {4'd10, 3'd2, 3'd1}: kernel_rom_out = 16'sd5462;
            {4'd10, 3'd2, 3'd2}: kernel_rom_out = 16'sd15937;
            {4'd10, 3'd2, 3'd3}: kernel_rom_out = -16'sd7178;
            {4'd10, 3'd2, 3'd4}: kernel_rom_out = 16'sd11876;
            {4'd10, 3'd2, 3'd5}: kernel_rom_out = -16'sd21097;
            {4'd10, 3'd2, 3'd6}: kernel_rom_out = 16'sd3226;
            {4'd10, 3'd2, 3'd7}: kernel_rom_out = -16'sd3346;
            {4'd10, 3'd3, 3'd0}: kernel_rom_out = -16'sd11902;
            {4'd10, 3'd3, 3'd1}: kernel_rom_out = -16'sd14876;
            {4'd10, 3'd3, 3'd2}: kernel_rom_out = -16'sd6159;
            {4'd10, 3'd3, 3'd3}: kernel_rom_out = 16'sd4114;
            {4'd10, 3'd3, 3'd4}: kernel_rom_out = -16'sd8012;
            {4'd10, 3'd3, 3'd5}: kernel_rom_out = -16'sd7623;
            {4'd10, 3'd3, 3'd6}: kernel_rom_out = -16'sd15508;
            {4'd10, 3'd3, 3'd7}: kernel_rom_out = -16'sd17119;
            {4'd10, 3'd4, 3'd0}: kernel_rom_out = -16'sd11902;
            {4'd10, 3'd4, 3'd1}: kernel_rom_out = 16'sd14876;
            {4'd10, 3'd4, 3'd2}: kernel_rom_out = -16'sd6159;
            {4'd10, 3'd4, 3'd3}: kernel_rom_out = -16'sd4114;
            {4'd10, 3'd4, 3'd4}: kernel_rom_out = -16'sd8012;
            {4'd10, 3'd4, 3'd5}: kernel_rom_out = 16'sd7623;
            {4'd10, 3'd4, 3'd6}: kernel_rom_out = 16'sd15508;
            {4'd10, 3'd4, 3'd7}: kernel_rom_out = -16'sd17119;
            {4'd10, 3'd5, 3'd0}: kernel_rom_out = -16'sd11428;
            {4'd10, 3'd5, 3'd1}: kernel_rom_out = -16'sd5462;
            {4'd10, 3'd5, 3'd2}: kernel_rom_out = 16'sd15937;
            {4'd10, 3'd5, 3'd3}: kernel_rom_out = 16'sd7178;
            {4'd10, 3'd5, 3'd4}: kernel_rom_out = 16'sd11876;
            {4'd10, 3'd5, 3'd5}: kernel_rom_out = 16'sd21097;
            {4'd10, 3'd5, 3'd6}: kernel_rom_out = -16'sd3226;
            {4'd10, 3'd5, 3'd7}: kernel_rom_out = -16'sd3346;
            {4'd10, 3'd6, 3'd0}: kernel_rom_out = -16'sd11768;
            {4'd10, 3'd6, 3'd1}: kernel_rom_out = -16'sd6617;
            {4'd10, 3'd6, 3'd2}: kernel_rom_out = -16'sd14607;
            {4'd10, 3'd6, 3'd3}: kernel_rom_out = 16'sd16824;
            {4'd10, 3'd6, 3'd4}: kernel_rom_out = 16'sd10658;
            {4'd10, 3'd6, 3'd5}: kernel_rom_out = -16'sd5380;
            {4'd10, 3'd6, 3'd6}: kernel_rom_out = 16'sd13456;
            {4'd10, 3'd6, 3'd7}: kernel_rom_out = 16'sd8449;
            {4'd10, 3'd7, 3'd0}: kernel_rom_out = -16'sd11229;
            {4'd10, 3'd7, 3'd1}: kernel_rom_out = 16'sd15554;
            {4'd10, 3'd7, 3'd2}: kernel_rom_out = 16'sd5617;
            {4'd10, 3'd7, 3'd3}: kernel_rom_out = 16'sd13614;
            {4'd10, 3'd7, 3'd4}: kernel_rom_out = -16'sd14765;
            {4'd10, 3'd7, 3'd5}: kernel_rom_out = -16'sd2171;
            {4'd10, 3'd7, 3'd6}: kernel_rom_out = -16'sd10240;
            {4'd10, 3'd7, 3'd7}: kernel_rom_out = 16'sd12696;

            // MODE 11: RFT-ENTROPY (unitarity: 1.80e-15)
            {4'd11, 3'd0, 3'd0}: kernel_rom_out = -16'sd14051;
            {4'd11, 3'd0, 3'd1}: kernel_rom_out = -16'sd2494;
            {4'd11, 3'd0, 3'd2}: kernel_rom_out = 16'sd18787;
            {4'd11, 3'd0, 3'd3}: kernel_rom_out = -16'sd9991;
            {4'd11, 3'd0, 3'd4}: kernel_rom_out = -16'sd4227;
            {4'd11, 3'd0, 3'd5}: kernel_rom_out = -16'sd14890;
            {4'd11, 3'd0, 3'd6}: kernel_rom_out = 16'sd11475;
            {4'd11, 3'd0, 3'd7}: kernel_rom_out = -16'sd6781;
            {4'd11, 3'd1, 3'd0}: kernel_rom_out = -16'sd1723;
            {4'd11, 3'd1, 3'd1}: kernel_rom_out = -16'sd16243;
            {4'd11, 3'd1, 3'd2}: kernel_rom_out = 16'sd4200;
            {4'd11, 3'd1, 3'd3}: kernel_rom_out = 16'sd20030;
            {4'd11, 3'd1, 3'd4}: kernel_rom_out = -16'sd1295;
            {4'd11, 3'd1, 3'd5}: kernel_rom_out = -16'sd11445;
            {4'd11, 3'd1, 3'd6}: kernel_rom_out = -16'sd14446;
            {4'd11, 3'd1, 3'd7}: kernel_rom_out = -16'sd6833;
            {4'd11, 3'd2, 3'd0}: kernel_rom_out = 16'sd14915;
            {4'd11, 3'd2, 3'd1}: kernel_rom_out = -16'sd6872;
            {4'd11, 3'd2, 3'd2}: kernel_rom_out = -16'sd12760;
            {4'd11, 3'd2, 3'd3}: kernel_rom_out = -16'sd3770;
            {4'd11, 3'd2, 3'd4}: kernel_rom_out = -16'sd15825;
            {4'd11, 3'd2, 3'd5}: kernel_rom_out = -16'sd7052;
            {4'd11, 3'd2, 3'd6}: kernel_rom_out = 16'sd10854;
            {4'd11, 3'd2, 3'd7}: kernel_rom_out = -16'sd14456;
            {4'd11, 3'd3, 3'd0}: kernel_rom_out = 16'sd10675;
            {4'd11, 3'd3, 3'd1}: kernel_rom_out = 16'sd14818;
            {4'd11, 3'd3, 3'd2}: kernel_rom_out = 16'sd1849;
            {4'd11, 3'd3, 3'd3}: kernel_rom_out = -16'sd4649;
            {4'd11, 3'd3, 3'd4}: kernel_rom_out = 16'sd16336;
            {4'd11, 3'd3, 3'd5}: kernel_rom_out = -16'sd11593;
            {4'd11, 3'd3, 3'd6}: kernel_rom_out = -16'sd8869;
            {4'd11, 3'd3, 3'd7}: kernel_rom_out = -16'sd15336;
            {4'd11, 3'd4, 3'd0}: kernel_rom_out = -16'sd10675;
            {4'd11, 3'd4, 3'd1}: kernel_rom_out = 16'sd14818;
            {4'd11, 3'd4, 3'd2}: kernel_rom_out = 16'sd1849;
            {4'd11, 3'd4, 3'd3}: kernel_rom_out = 16'sd4649;
            {4'd11, 3'd4, 3'd4}: kernel_rom_out = -16'sd16336;
            {4'd11, 3'd4, 3'd5}: kernel_rom_out = 16'sd11593;
            {4'd11, 3'd4, 3'd6}: kernel_rom_out = -16'sd8869;
            {4'd11, 3'd4, 3'd7}: kernel_rom_out = -16'sd15336;
            {4'd11, 3'd5, 3'd0}: kernel_rom_out = -16'sd14915;
            {4'd11, 3'd5, 3'd1}: kernel_rom_out = -16'sd6872;
            {4'd11, 3'd5, 3'd2}: kernel_rom_out = -16'sd12760;
            {4'd11, 3'd5, 3'd3}: kernel_rom_out = 16'sd3770;
            {4'd11, 3'd5, 3'd4}: kernel_rom_out = 16'sd15825;
            {4'd11, 3'd5, 3'd5}: kernel_rom_out = 16'sd7052;
            {4'd11, 3'd5, 3'd6}: kernel_rom_out = 16'sd10854;
            {4'd11, 3'd5, 3'd7}: kernel_rom_out = -16'sd14456;
            {4'd11, 3'd6, 3'd0}: kernel_rom_out = 16'sd1723;
            {4'd11, 3'd6, 3'd1}: kernel_rom_out = -16'sd16243;
            {4'd11, 3'd6, 3'd2}: kernel_rom_out = 16'sd4200;
            {4'd11, 3'd6, 3'd3}: kernel_rom_out = -16'sd20030;
            {4'd11, 3'd6, 3'd4}: kernel_rom_out = 16'sd1295;
            {4'd11, 3'd6, 3'd5}: kernel_rom_out = 16'sd11445;
            {4'd11, 3'd6, 3'd6}: kernel_rom_out = -16'sd14446;
            {4'd11, 3'd6, 3'd7}: kernel_rom_out = -16'sd6833;
            {4'd11, 3'd7, 3'd0}: kernel_rom_out = 16'sd14051;
            {4'd11, 3'd7, 3'd1}: kernel_rom_out = -16'sd2494;
            {4'd11, 3'd7, 3'd2}: kernel_rom_out = 16'sd18787;
            {4'd11, 3'd7, 3'd3}: kernel_rom_out = 16'sd9991;
            {4'd11, 3'd7, 3'd4}: kernel_rom_out = 16'sd4227;
            {4'd11, 3'd7, 3'd5}: kernel_rom_out = 16'sd14890;
            {4'd11, 3'd7, 3'd6}: kernel_rom_out = 16'sd11475;
            {4'd11, 3'd7, 3'd7}: kernel_rom_out = -16'sd6781;

            default: kernel_rom_out = 16'sd11585;
        endcase
    end

    // Clock/reset
    always @(posedge WF_CLK) begin
        if (reset_counter < 8'd10)
            reset_counter <= reset_counter + 1'b1;
    end
    
    always @(posedge WF_CLK) begin
        if (reset) begin
            button_debounce <= 20'h00000;
            button_stable <= 1'b0;
            button_prev <= 1'b0;
        end else begin
            button_debounce <= {button_debounce[18:0], ~WF_BUTTON};
            button_stable <= &button_debounce[19:16];
            button_prev <= button_stable;
        end
    end
    
    always @(posedge WF_CLK) begin
        if (reset) begin
            current_mode <= MODE_RFT_GOLDEN;
            auto_cycle_counter <= 24'h000000;
        end else begin
            auto_cycle_counter <= auto_cycle_counter + 1'b1;
            if (button_edge || auto_cycle_trigger) begin
                current_mode <= current_mode + 1'b1;
                auto_cycle_counter <= 24'h000000;
            end
        end
    end
    
    always @(posedge WF_CLK) begin
        if (reset)
            cyc_cnt <= 8'h00;
        else
            cyc_cnt <= cyc_cnt + 1'b1;
    end

    // Input data (ramp pattern)
    always @(posedge WF_CLK) begin
        if (reset) begin
            for (i = 0; i < 8; i = i + 1)
                sample[i] <= 16'h0000;
            valid <= 1'b0;
        end
        else if (start && !valid) begin
            sample[0] <= 16'h0000;
            sample[1] <= 16'h1000;
            sample[2] <= 16'h2000;
            sample[3] <= 16'h3000;
            sample[4] <= 16'h4000;
            sample[5] <= 16'h5000;
            sample[6] <= 16'h6000;
            sample[7] <= 16'h7000;
            valid <= 1'b1;
        end
    end

    // State machine
    always @(posedge WF_CLK) begin
        if (reset) begin
            state <= STATE_IDLE;
            k_index <= 3'b000;
            n_index <= 3'b000;
        end
        else begin
            case (state)
                STATE_IDLE: begin
                    if (start) begin
                        k_index <= 3'b000;
                        n_index <= 3'b000;
                        state <= STATE_COMPUTE;
                    end
                end
                
                STATE_COMPUTE: begin
                    if (n_index == 3'b111) begin
                        if (k_index == 3'b111)
                            state <= STATE_DONE;
                        else begin
                            k_index <= k_index + 1'b1;
                            n_index <= 3'b000;
                        end
                    end
                    else
                        n_index <= n_index + 1'b1;
                end
                
                STATE_DONE: state <= STATE_IDLE;
                
                default: state <= STATE_IDLE;
            endcase
        end
    end

    // Pipeline register for kernel
    always @(posedge WF_CLK) begin
        kernel_reg <= kernel_rom_out;
    end

    // Accumulator
    always @(posedge WF_CLK) begin
        if (reset || state == STATE_IDLE)
            acc <= 32'sh00000000;
        else if (is_computing) begin
            if (n_index == 3'b000)
                acc <= mult_out;
            else
                acc <= acc + mult_out;
        end
    end

    // Result storage
    always @(posedge WF_CLK) begin
        if (reset) begin
            for (i = 0; i < 8; i = i + 1)
                rft_out[i] <= 32'sh00000000;
        end
        else if (save_result)
            rft_out[k_index] <= acc;
    end

    // Magnitude
    wire [31:0] amplitude [0:7];
    genvar g;
    generate
        for (g = 0; g < 8; g = g + 1) begin : mag_calc
            assign amplitude[g] = rft_out[g][31] ? -rft_out[g] : rft_out[g];
        end
    endgenerate

    // LED output
    always @(posedge WF_CLK) begin
        if (reset)
            led_output <= 8'h00;
        else if (is_done) begin
            led_output[0] <= (amplitude[0][30:23] > 8'd32);
            led_output[1] <= (amplitude[1][30:23] > 8'd16);
            led_output[2] <= (amplitude[2][30:23] > 8'd8);
            led_output[3] <= (amplitude[3][30:23] > 8'd8);
            led_output[4] <= (amplitude[4][30:23] > 8'd8);
            led_output[5] <= (amplitude[5][30:23] > 8'd8);
            led_output[6] <= (amplitude[6][30:23] > 8'd16);
            led_output[7] <= (amplitude[7][30:23] > 8'd32);
        end
        else
            led_output <= {4'b0000, current_mode};
    end
    
    assign WF_LED = led_output;

endmodule
